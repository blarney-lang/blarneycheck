module top (
  input wire clock,
  input wire reset
  );
  // Declarations
  //////////////////////////////////////////////////////////////////////////////
  wire [0:0] v_0_0;
  wire [0:0] v_1_0;
  wire [0:0] v_2_0;
  reg [2:0] v_3_0 = 3'h0;
  wire [0:0] v_4_0;
  wire [0:0] v_5_0;
  wire [0:0] v_6_0;
  wire [0:0] v_7_0;
  reg [0:0] v_8_0 = 1'h1;
  wire [0:0] v_9_0;
  wire [0:0] v_10_0;
  wire [0:0] v_11_0;
  wire [0:0] v_12_0;
  wire [0:0] v_13_0;
  wire [0:0] v_14_0;
  wire [0:0] v_15_0;
  reg [0:0] v_16_0 = 1'h0;
  wire [0:0] v_17_0;
  wire [0:0] v_18_0;
  wire [0:0] v_19_0;
  wire [0:0] v_20_0;
  reg [0:0] v_21_0 = 1'h0;
  wire [0:0] v_22_0;
  wire [0:0] v_23_0;
  wire [0:0] v_24_0;
  wire [0:0] v_25_0;
  wire [0:0] v_26_0;
  wire [0:0] v_27_0;
  wire [0:0] v_28_0;
  wire [0:0] v_29_0;
  wire [0:0] v_30_0;
  wire [0:0] v_31_0;
  wire [0:0] v_32_0;
  wire [4:0] v_33_0;
   wire [4:0] v_34_0;
  wire [7:0] v_35_0;
  wire [7:0] v_36_0;
  wire [7:0] v_37_0;
  reg [7:0] v_38_0 = 8'h0;
  wire [0:0] v_39_0;
  wire [0:0] v_40_0;
  wire [0:0] v_41_0;
  wire [0:0] v_42_0;
  wire [0:0] v_43_0;
  wire [7:0] v_44_0;
  wire [7:0] v_45_0;
  wire [7:0] v_46_0;
  wire [7:0] v_47_0;
  wire [7:0] v_48_0;
  wire [7:0] v_49_0;
  wire [7:0] v_50_0;
  wire [7:0] v_51_0;
  wire [7:0] v_52_0;
  wire [7:0] v_53_0;
  wire [7:0] v_54_0;
  wire [7:0] v_55_0;
  wire [7:0] v_56_0;
  wire [0:0] v_57_0;
  wire [0:0] v_58_0;
  wire [0:0] v_59_0;
  wire [0:0] v_60_0;
  wire [7:0] v_61_0;
  wire [7:0] v_62_0;
  wire [7:0] v_63_0;
  wire [4:0] v_64_0;
  wire [4:0] v_65_0;
  wire [0:0] v_66_0;
  wire [0:0] v_67_0;
  wire [4:0] v_68_0;
  wire [4:0] v_69_0;
  wire [4:0] v_70_0;
  wire [4:0] v_71_0;
  wire [0:0] v_72_0;
  wire [0:0] v_73_0;
  wire [0:0] v_74_0;
  wire [0:0] v_75_0;
  wire [0:0] v_76_0;
  wire [0:0] v_77_0;
  wire [0:0] v_78_0;
  wire [0:0] v_79_0;
  wire [0:0] v_80_0;
  wire [0:0] v_81_0;
  wire [0:0] v_82_0;
  wire [0:0] v_83_0;
  wire [0:0] v_84_0;
  wire [0:0] v_85_0;
  wire [0:0] v_86_0;
  wire [0:0] v_87_0;
  wire [0:0] v_88_0;
  wire [0:0] v_89_0;
  wire [0:0] v_90_0;
  wire [0:0] v_91_0;
  wire [0:0] v_92_0;
  wire [0:0] v_93_0;
  wire [0:0] v_94_0;
  wire [0:0] v_95_0;
  wire [0:0] v_96_0;
  wire [0:0] v_97_0;
  wire [0:0] v_98_0;
  wire [0:0] v_99_0;
  wire [0:0] v_100_0;
  wire [0:0] v_101_0;
  wire [0:0] v_102_0;
  wire [0:0] v_103_0;
  wire [0:0] v_104_0;
  wire [0:0] v_105_0;
  wire [0:0] v_106_0;
  wire [2:0] v_107_0;
  wire [2:0] v_108_0;
  wire [2:0] v_109_0;
  wire [2:0] v_110_0;
  wire [0:0] v_113_0;
  reg [0:0] v_114_0 = 1'h0;
  wire [0:0] v_115_0;
  // Instances
  //////////////////////////////////////////////////////////////////////////////
  assign v_0_0 = v_1_0 & v_7_0;
  assign v_1_0 = ~(v_2_0);
  assign v_2_0 = v_3_0 != 3'h9;
  assign v_4_0 = v_5_0 | v_105_0;
  assign v_5_0 = v_6_0 & v_104_0;
  assign v_6_0 = v_7_0 & v_103_0;
  assign v_7_0 = 1'h1 & v_8_0;
  assign v_9_0 = v_10_0 | v_95_0;
  assign v_10_0 = v_11_0 & v_21_0;
  assign v_11_0 = v_12_0 & v_94_0;
  assign v_12_0 = v_13_0 & v_15_0;
  assign v_13_0 = 1'h1 & v_14_0;
  assign v_14_0 = ~(v_8_0);
  assign v_15_0 = ~(v_16_0);
  assign v_17_0 = v_18_0 | v_42_0;
  assign v_18_0 = v_19_0 & v_90_0;
  assign v_19_0 = v_20_0 & v_21_0;
  assign v_20_0 = v_13_0 & v_16_0;
  assign v_22_0 = v_23_0 | v_26_0;
  assign v_23_0 = v_24_0 | v_10_0;
  assign v_24_0 = v_20_0 & v_25_0;
  assign v_25_0 = ~(v_21_0);
  assign v_26_0 = v_27_0 | v_29_0;
  assign v_27_0 = v_11_0 & v_28_0;
  assign v_28_0 = ~(v_21_0);
  assign v_29_0 = v_30_0 | v_18_0;
  assign v_30_0 = v_31_0 & v_79_0;
  assign v_31_0 = v_19_0 & v_32_0;
  assign v_32_0 = 5'h0 <= v_33_0;
  assign v_33_0 = v_34_0 + 5'h1;
  BlockRAM# (
      .INIT_FILE("UNUSED"),
      .ADDR_WIDTH(8),
      .DATA_WIDTH(5)
    ) ram34 (
      .CLK(clock),
      .DI(v_64_0),
      .ADDR(v_35_0),
      .WE(v_72_0),
      .DO(v_34_0)
    );
  assign v_35_0 = v_36_0 | v_55_0;
  assign v_36_0 = v_37_0 | v_54_0;
  assign v_37_0 = v_24_0 ? v_38_0 : 8'h0;
  assign v_39_0 = v_40_0 | v_41_0;
  assign v_40_0 = v_30_0 | v_18_0;
  assign v_41_0 = v_42_0 | v_10_0;
  assign v_42_0 = v_12_0 & v_43_0;
  assign v_43_0 = 8'h0 < v_38_0;
  assign v_44_0 = v_45_0 | v_49_0;
  assign v_45_0 = v_46_0 | v_48_0;
  assign v_46_0 = v_30_0 ? v_47_0 : 8'h0;
  assign v_47_0 = v_38_0 - 8'h1;
  assign v_48_0 = v_18_0 ? 8'h0 : 8'h0;
  assign v_49_0 = v_50_0 | v_52_0;
  assign v_50_0 = v_42_0 ? v_51_0 : 8'h0;
  assign v_51_0 = v_38_0 - 8'h1;
  assign v_52_0 = v_10_0 ? v_53_0 : 8'h0;
  assign v_53_0 = v_38_0 + 8'h1;
  assign v_54_0 = v_27_0 ? v_38_0 : 8'h0;
  assign v_55_0 = v_56_0 | v_61_0;
  assign v_56_0 = v_57_0 ? 8'bxxxxxxxx : 8'h0;
  assign v_57_0 = ~(v_58_0);
  assign v_58_0 = v_59_0 | v_60_0;
  assign v_59_0 = v_30_0 | v_18_0;
  assign v_60_0 = v_24_0 | v_27_0;
  assign v_61_0 = v_62_0 | v_63_0;
  assign v_62_0 = v_30_0 ? v_38_0 : 8'h0;
  assign v_63_0 = v_18_0 ? v_38_0 : 8'h0;
  assign v_64_0 = v_65_0 | v_68_0;
  assign v_65_0 = v_66_0 ? 5'bxxxxx : 5'h0;
  assign v_66_0 = ~(v_67_0);
  assign v_67_0 = v_30_0 | v_18_0;
  assign v_68_0 = v_69_0 | v_70_0;
  assign v_69_0 = v_30_0 ? 5'h0 : 5'h0;
  assign v_70_0 = v_18_0 ? v_71_0 : 5'h0;
  assign v_71_0 = v_34_0 + 5'h1;
  assign v_72_0 = v_73_0 | v_76_0;
  assign v_73_0 = v_74_0 ? 1'h0 : 1'h0;
  assign v_74_0 = ~(v_75_0);
  assign v_75_0 = v_30_0 | v_18_0;
  assign v_76_0 = v_77_0 | v_78_0;
  assign v_77_0 = v_30_0 ? 1'h1 : 1'h0;
  assign v_78_0 = v_18_0 ? 1'h1 : 1'h0;
  assign v_79_0 = ~(v_80_0);
  assign v_80_0 = v_38_0 == 8'h0;
  assign v_81_0 = v_82_0 | v_85_0;
  assign v_82_0 = v_83_0 | v_84_0;
  assign v_83_0 = v_24_0 ? 1'h1 : 1'h0;
  assign v_84_0 = v_10_0 ? 1'h0 : 1'h0;
  assign v_85_0 = v_86_0 | v_87_0;
  assign v_86_0 = v_27_0 ? 1'h1 : 1'h0;
  assign v_87_0 = v_88_0 | v_89_0;
  assign v_88_0 = v_30_0 ? 1'h0 : 1'h0;
  assign v_89_0 = v_18_0 ? 1'h0 : 1'h0;
  assign v_90_0 = ~(v_32_0);
  assign v_91_0 = v_92_0 | v_93_0;
  assign v_92_0 = v_18_0 ? 1'h0 : 1'h0;
  assign v_93_0 = v_42_0 ? 1'h1 : 1'h0;
  assign v_94_0 = ~(v_43_0);
  assign v_95_0 = v_7_0 | v_18_0;
  assign v_96_0 = v_97_0 | v_98_0;
  assign v_97_0 = v_10_0 ? 1'h1 : 1'h0;
  assign v_98_0 = v_99_0 | v_102_0;
  assign v_99_0 = v_7_0 ? v_100_0 : 1'h0;
  assign v_100_0 = v_101_0 & 1'h1;
  assign v_101_0 = v_3_0 != 3'h7;
  assign v_102_0 = v_18_0 ? 1'h1 : 1'h0;
  assign v_103_0 = v_3_0 != 3'h7;
  assign v_104_0 = ~(1'h1);
  assign v_105_0 = v_7_0 & v_106_0;
  assign v_106_0 = ~(v_103_0);
  assign v_107_0 = v_108_0 | v_109_0;
  assign v_108_0 = v_5_0 ? 3'h0 : 3'h0;
  assign v_109_0 = v_105_0 ? v_110_0 : 3'h0;
  assign v_110_0 = v_3_0 + 3'h1;
  assign v_113_0 = v_114_0 & 1'h1;
  assign v_115_0 = v_31_0 & v_80_0;
  // Always block
  //////////////////////////////////////////////////////////////////////////////
  always @(posedge clock) begin
    if (reset) begin
      v_3_0 <= 3'h0;
      v_8_0 <= 1'h1;
      v_16_0 <= 1'h0;
      v_21_0 <= 1'h0;
      v_38_0 <= 8'h0;
      v_114_0 <= 1'h0;
    end else begin
      if (v_4_0 == 1) v_3_0 <= v_107_0;
      if (v_9_0 == 1) v_8_0 <= v_96_0;
      if (v_17_0 == 1) v_16_0 <= v_91_0;
      if (v_22_0 == 1) v_21_0 <= v_81_0;
      if (v_39_0 == 1) v_38_0 <= v_44_0;
      if (v_0_0 == 1) $write (
        "Test",
        "=",
        v_3_0,
        ", "
      );
      if (v_0_0 == 1) $write (
        "Failed the test.",
        "\n"
      );
      if (v_115_0 == 1) v_114_0 <= 1'h1;
      if (v_113_0 == 1) $finish;
      if (v_0_0 == 1) $finish;
    end
  end
endmodule