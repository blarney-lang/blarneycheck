module Top
  (input wire clock,
   input wire reset,
   input wire [0:0] in_canPeek,
   input wire [0:0] out_consume_en,
   input wire [7:0] in_peek,
   output wire [0:0] in_consume_en,
   output wire [0:0] out_canPeek,
   output wire [7:0] out_peek);
  // Declarations
  //////////////////////////////////////////////////////////////////////////////
  wire [0:0] v_1_0;
  wire [0:0] v_2_0;
  reg [0:0] v_3_0 = 1'h0;
  wire [0:0] v_4_0;
  wire [0:0] v_5_0;
  wire [0:0] v_6_0;
  wire [0:0] v_7_0;
  wire [0:0] v_8_0;
  wire [0:0] v_9_0;
  wire [15:0] v_10_0;
  wire [0:0] v_11_0;
  reg [15:0] v_12_0 = 16'h0;
  wire [0:0] v_13_0;
  wire [0:0] v_14_0;
  wire [0:0] v_15_0;
  wire [0:0] v_16_0;
  wire [0:0] v_17_0;
  reg [0:0] v_18_0 = 1'h0;
  wire [0:0] v_19_0;
  wire [0:0] v_20_0;
  wire [0:0] v_21_0;
  wire [0:0] v_22_0;
  reg [9:0] v_23_0 = 10'h0;
  wire [0:0] v_24_0;
  wire [0:0] v_25_0;
  wire [0:0] v_26_0;
  wire [0:0] v_27_0;
  wire [0:0] v_28_0;
  wire [0:0] v_29_0;
  wire [0:0] v_30_0;
  wire [0:0] v_31_0;
  wire [0:0] v_32_0;
  wire [0:0] v_33_0;
  reg [0:0] v_34_0 = 1'h1;
  wire [0:0] v_35_0;
  wire [0:0] v_36_0;
  wire [0:0] v_37_0;
  wire [0:0] v_38_0;
  wire [0:0] v_39_0;
  reg [0:0] v_40_0 = 1'h1;
  wire [0:0] v_41_0;
  wire [0:0] v_42_0;
  wire [0:0] v_43_0;
  wire [0:0] v_44_0;
  wire [0:0] v_45_0;
  wire [0:0] v_46_0;
  wire [0:0] v_47_0;
  wire [0:0] v_48_0;
  wire [0:0] v_49_0;
  wire [2:0] v_50_0;
  wire [0:0] v_51_0;
  reg [15:0] v_52_0 = 16'h0;
  wire [15:0] v_53_0;
  reg [2:0] v_54_0 = 3'h0;
  wire [0:0] v_55_0;
  wire [0:0] v_56_0;
  wire [0:0] v_57_0;
  reg [0:0] v_58_0 = 1'h0;
  wire [0:0] v_59_0;
  reg [0:0] v_60_0 = 1'h0;
  wire [0:0] v_61_0;
  wire [0:0] v_62_0;
  wire [0:0] _act_63_0;
  wire [0:0] v_64_0;
  wire [0:0] v_65_0;
  wire [0:0] v_66_0;
  reg [0:0] v_67_0 = 1'h1;
  wire [0:0] v_68_0;
  wire [0:0] v_69_0;
  wire [0:0] v_70_0;
  wire [4:0] v_71_0;
  wire [0:0] v_72_0;
  wire [0:0] v_73_0;
  wire [0:0] v_74_0;
  wire [0:0] v_75_0;
  wire [4:0] v_76_0;
  reg [4:0] v_77_0 = 5'h0;
  reg [4:0] v_78_0 = 5'h0;
  wire [0:0] _act_79_0;
  wire [0:0] _act_80_0;
  wire [0:0] v_81_0;
  wire [0:0] v_82_0;
  wire [0:0] v_83_0;
  wire [0:0] v_84_0;
  wire [0:0] v_85_0;
  wire [0:0] v_86_0;
  wire [0:0] v_87_0;
  wire [0:0] v_88_0;
  wire [0:0] v_89_0;
  wire [0:0] v_90_0;
  reg [0:0] v_91_0 = 1'h0;
  wire [0:0] v_92_0;
  wire [0:0] v_93_0;
  wire [0:0] v_94_0;
  wire [0:0] v_95_0;
  wire [15:0] v_96_0;
  reg [15:0] v_97_0 = 16'h0;
  wire [0:0] v_98_0;
  wire [0:0] v_99_0;
  wire [0:0] v_100_0;
  wire [0:0] v_101_0;
  wire [0:0] v_102_0;
  wire [0:0] v_103_0;
  wire [0:0] v_104_0;
  wire [15:0] v_105_0;
  wire [15:0] v_106_0;
  wire [15:0] v_107_0;
  wire [15:0] v_108_0;
  wire [15:0] v_109_0;
  wire [15:0] v_110_0;
  wire [15:0] v_111_0;
  wire [15:0] v_112_0;
  wire [15:0] v_113_0;
  wire [0:0] v_114_0;
  wire [0:0] v_115_0;
  wire [0:0] v_116_0;
  wire [0:0] v_117_0;
  wire [0:0] v_118_0;
  wire [0:0] v_119_0;
  wire [0:0] v_120_0;
  wire [0:0] v_121_0;
  wire [0:0] v_122_0;
  wire [0:0] v_123_0;
  wire [0:0] v_124_0;
  wire [0:0] v_125_0;
  wire [0:0] v_126_0;
  wire [0:0] v_127_0;
  wire [0:0] v_128_0;
  wire [0:0] v_129_0;
  wire [0:0] v_130_0;
  wire [0:0] v_131_0;
  wire [0:0] v_132_0;
  wire [0:0] v_133_0;
  wire [0:0] v_134_0;
  wire [0:0] v_135_0;
  wire [0:0] v_136_0;
  wire [0:0] v_137_0;
  wire [0:0] v_138_0;
  wire [0:0] v_139_0;
  wire [0:0] v_140_0;
  wire [0:0] v_141_0;
  wire [0:0] v_142_0;
  wire [0:0] v_143_0;
  wire [0:0] v_144_0;
  wire [0:0] v_145_0;
  wire [0:0] v_146_0;
  wire [0:0] v_147_0;
  wire [0:0] v_148_0;
  wire [0:0] v_149_0;
  wire [0:0] v_150_0;
  wire [0:0] v_151_0;
  wire [0:0] v_152_0;
  wire [0:0] v_153_0;
  wire [0:0] v_154_0;
  wire [0:0] v_155_0;
  wire [0:0] v_156_0;
  wire [0:0] v_157_0;
  wire [0:0] v_158_0;
  wire [0:0] v_159_0;
  wire [0:0] v_160_0;
  wire [0:0] v_161_0;
  wire [4:0] v_162_0;
  wire [0:0] v_163_0;
  wire [0:0] v_164_0;
  wire [0:0] v_165_0;
  wire [0:0] v_166_0;
  wire [0:0] v_167_0;
  wire [0:0] v_168_0;
  wire [0:0] v_169_0;
  wire [0:0] v_170_0;
  wire [0:0] v_171_0;
  wire [0:0] v_172_0;
  wire [0:0] v_173_0;
  wire [0:0] v_174_0;
  wire [0:0] v_175_0;
  wire [0:0] v_176_0;
  wire [0:0] v_177_0;
  wire [0:0] v_178_0;
  wire [0:0] v_179_0;
  wire [0:0] v_180_0;
  wire [0:0] v_181_0;
  wire [0:0] v_182_0;
  wire [0:0] v_183_0;
  wire [0:0] v_184_0;
  wire [0:0] v_185_0;
  wire [0:0] v_186_0;
  wire [0:0] v_187_0;
  wire [0:0] v_188_0;
  wire [0:0] v_189_0;
  wire [2:0] v_190_0;
  reg [2:0] v_191_0 = 3'h0;
  wire [0:0] v_192_0;
  wire [0:0] v_193_0;
  wire [0:0] v_194_0;
  wire [0:0] v_195_0;
  wire [0:0] v_196_0;
  wire [0:0] v_197_0;
  wire [0:0] v_198_0;
  wire [0:0] v_199_0;
  wire [2:0] v_200_0;
  wire [2:0] v_201_0;
  wire [2:0] v_202_0;
  wire [0:0] v_203_0;
  wire [0:0] v_204_0;
  reg [0:0] v_205_0 = 1'h0;
  reg [0:0] v_206_0 = 1'h0;
  wire [0:0] v_207_0;
  reg [4:0] v_208_0 = 5'h0;
  wire [4:0] v_209_0;
  wire [4:0] v_210_0;
  wire [4:0] v_211_0;
  wire [0:0] v_212_0;
  reg [4:0] v_213_0 = 5'h0;
  wire [4:0] v_214_0;
  wire [4:0] v_215_0;
  wire [4:0] v_216_0;
  wire [0:0] v_217_0;
  reg [2:0] v_218_0 = 3'h0;
  wire [2:0] v_219_0;
  wire [2:0] v_220_0;
  wire [2:0] v_221_0;
  wire [2:0] v_222_0;
  wire [2:0] v_223_0;
  wire [2:0] v_224_0;
  wire [2:0] v_225_0;
  wire [2:0] v_226_0;
  wire [2:0] v_227_0;
  wire [2:0] v_228_0;
  wire [2:0] v_229_0;
  wire [2:0] v_230_0;
  wire [2:0] v_231_0;
  wire [2:0] v_232_0;
  wire [0:0] v_233_0;
  wire [2:0] v_234_0;
  wire [2:0] v_235_0;
  wire [2:0] v_236_0;
  wire [2:0] v_237_0;
  wire [2:0] v_238_0;
  wire [2:0] v_239_0;
  wire [2:0] v_240_0;
  wire [2:0] v_241_0;
  wire [2:0] v_242_0;
  wire [2:0] v_243_0;
  wire [2:0] v_244_0;
  wire [2:0] v_245_0;
  wire [2:0] v_246_0;
  wire [0:0] v_247_0;
  wire [2:0] v_248_0;
  wire [2:0] v_248_1;
  wire [4:0] v_249_0;
  wire [4:0] v_250_0;
  wire [4:0] v_251_0;
  wire [0:0] v_252_0;
  wire [2:0] v_253_0;
  wire [0:0] v_254_0;
  wire [0:0] v_255_0;
  wire [0:0] v_256_0;
  wire [4:0] v_257_0;
  wire [4:0] v_258_0;
  wire [4:0] v_259_0;
  wire [0:0] v_260_0;
  wire [2:0] v_261_0;
  wire [2:0] v_262_0;
  wire [2:0] v_263_0;
  wire [0:0] v_264_0;
  wire [0:0] v_265_0;
  wire [0:0] v_266_0;
  wire [0:0] v_267_0;
  wire [0:0] v_268_0;
  wire [2:0] v_269_0;
  wire [0:0] v_270_0;
  reg [2:0] v_271_0 = 3'h0;
  wire [0:0] v_272_0;
  wire [0:0] v_273_0;
  wire [0:0] v_274_0;
  wire [0:0] v_275_0;
  wire [0:0] v_276_0;
  wire [0:0] v_277_0;
  wire [0:0] v_278_0;
  wire [0:0] v_279_0;
  wire [0:0] v_280_0;
  wire [0:0] v_281_0;
  wire [0:0] v_282_0;
  wire [0:0] v_283_0;
  wire [0:0] v_284_0;
  wire [0:0] v_285_0;
  wire [0:0] v_286_0;
  wire [0:0] v_287_0;
  wire [0:0] v_288_0;
  wire [0:0] v_289_0;
  wire [0:0] v_290_0;
  wire [0:0] v_291_0;
  wire [0:0] v_292_0;
  wire [0:0] v_293_0;
  wire [0:0] v_294_0;
  wire [0:0] v_295_0;
  wire [0:0] v_296_0;
  wire [0:0] v_297_0;
  wire [0:0] v_298_0;
  wire [0:0] v_299_0;
  wire [0:0] v_300_0;
  wire [2:0] v_301_0;
  wire [2:0] v_302_0;
  wire [2:0] v_303_0;
  wire [2:0] v_304_0;
  wire [2:0] v_305_0;
  wire [2:0] v_306_0;
  wire [2:0] v_307_0;
  wire [2:0] v_308_0;
  wire [2:0] v_309_0;
  wire [2:0] v_310_0;
  wire [2:0] v_311_0;
  wire [2:0] v_312_0;
  wire [2:0] v_313_0;
  wire [2:0] v_314_0;
  wire [2:0] v_315_0;
  wire [2:0] v_316_0;
  wire [2:0] v_317_0;
  wire [2:0] v_318_0;
  wire [2:0] v_319_0;
  wire [0:0] v_320_0;
  wire [0:0] v_321_0;
  wire [0:0] v_322_0;
  wire [0:0] v_323_0;
  wire [0:0] v_324_0;
  wire [0:0] v_325_0;
  wire [0:0] v_326_0;
  wire [0:0] v_327_0;
  wire [2:0] v_328_0;
  wire [0:0] v_329_0;
  reg [15:0] v_330_0 = 16'h0;
  wire [15:0] v_331_0;
  reg [2:0] v_332_0 = 3'h0;
  wire [0:0] v_333_0;
  wire [0:0] v_334_0;
  wire [0:0] v_335_0;
  reg [0:0] v_336_0 = 1'h0;
  wire [0:0] v_337_0;
  reg [0:0] v_338_0 = 1'h0;
  wire [0:0] v_339_0;
  wire [0:0] v_340_0;
  wire [0:0] _act_341_0;
  wire [0:0] v_342_0;
  wire [0:0] v_343_0;
  wire [0:0] v_344_0;
  reg [0:0] v_345_0 = 1'h1;
  wire [0:0] v_346_0;
  wire [0:0] v_347_0;
  wire [0:0] v_348_0;
  wire [4:0] v_349_0;
  wire [0:0] v_350_0;
  wire [0:0] v_351_0;
  wire [0:0] v_352_0;
  wire [0:0] v_353_0;
  wire [4:0] v_354_0;
  reg [4:0] v_355_0 = 5'h0;
  reg [4:0] v_356_0 = 5'h0;
  wire [0:0] _act_357_0;
  wire [0:0] _act_358_0;
  wire [0:0] v_359_0;
  wire [0:0] v_360_0;
  wire [0:0] v_361_0;
  wire [0:0] v_362_0;
  wire [0:0] v_363_0;
  wire [0:0] v_364_0;
  wire [0:0] v_365_0;
  wire [0:0] v_366_0;
  wire [0:0] v_367_0;
  wire [0:0] v_368_0;
  wire [0:0] v_369_0;
  wire [0:0] v_370_0;
  wire [0:0] v_371_0;
  wire [0:0] v_372_0;
  wire [0:0] v_373_0;
  wire [0:0] v_374_0;
  wire [0:0] v_375_0;
  wire [0:0] v_376_0;
  wire [0:0] v_377_0;
  wire [0:0] v_378_0;
  wire [0:0] v_379_0;
  wire [0:0] v_380_0;
  wire [0:0] v_381_0;
  wire [0:0] v_382_0;
  wire [0:0] v_383_0;
  wire [0:0] v_384_0;
  wire [0:0] v_385_0;
  wire [0:0] v_386_0;
  wire [0:0] v_387_0;
  wire [0:0] v_388_0;
  wire [0:0] v_389_0;
  wire [0:0] v_390_0;
  wire [0:0] v_391_0;
  wire [0:0] v_392_0;
  wire [0:0] v_393_0;
  wire [0:0] v_394_0;
  wire [0:0] v_395_0;
  wire [0:0] v_396_0;
  wire [0:0] v_397_0;
  wire [0:0] v_398_0;
  wire [0:0] v_399_0;
  wire [0:0] v_400_0;
  wire [0:0] v_401_0;
  wire [0:0] v_402_0;
  wire [0:0] v_403_0;
  wire [0:0] v_404_0;
  wire [4:0] v_405_0;
  wire [0:0] v_406_0;
  wire [0:0] v_407_0;
  wire [0:0] v_408_0;
  wire [0:0] v_409_0;
  wire [0:0] v_410_0;
  wire [0:0] v_411_0;
  wire [0:0] v_412_0;
  wire [0:0] v_413_0;
  wire [0:0] v_414_0;
  wire [0:0] v_415_0;
  wire [0:0] v_416_0;
  wire [0:0] v_417_0;
  wire [0:0] v_418_0;
  wire [0:0] v_419_0;
  wire [0:0] v_420_0;
  wire [0:0] v_421_0;
  wire [0:0] v_422_0;
  wire [0:0] v_423_0;
  wire [0:0] v_424_0;
  wire [0:0] v_425_0;
  wire [0:0] v_426_0;
  wire [0:0] v_427_0;
  wire [0:0] v_428_0;
  wire [0:0] v_429_0;
  wire [0:0] v_430_0;
  wire [0:0] v_431_0;
  wire [0:0] v_432_0;
  wire [2:0] v_433_0;
  reg [2:0] v_434_0 = 3'h0;
  wire [0:0] v_435_0;
  wire [0:0] v_436_0;
  wire [0:0] v_437_0;
  wire [0:0] v_438_0;
  wire [0:0] v_439_0;
  wire [0:0] v_440_0;
  wire [0:0] v_441_0;
  wire [0:0] v_442_0;
  wire [2:0] v_443_0;
  wire [2:0] v_444_0;
  wire [2:0] v_445_0;
  wire [0:0] v_446_0;
  wire [0:0] v_447_0;
  reg [0:0] v_448_0 = 1'h0;
  reg [0:0] v_449_0 = 1'h0;
  wire [0:0] v_450_0;
  reg [4:0] v_451_0 = 5'h0;
  wire [4:0] v_452_0;
  wire [4:0] v_453_0;
  wire [4:0] v_454_0;
  wire [0:0] v_455_0;
  reg [4:0] v_456_0 = 5'h0;
  wire [4:0] v_457_0;
  wire [4:0] v_458_0;
  wire [4:0] v_459_0;
  wire [0:0] v_460_0;
  reg [2:0] v_461_0 = 3'h0;
  wire [2:0] v_462_0;
  wire [2:0] v_463_0;
  wire [2:0] v_464_0;
  wire [2:0] v_465_0;
  wire [2:0] v_466_0;
  wire [2:0] v_467_0;
  wire [2:0] v_468_0;
  wire [2:0] v_469_0;
  wire [2:0] v_470_0;
  wire [2:0] v_471_0;
  wire [2:0] v_472_0;
  wire [2:0] v_473_0;
  wire [2:0] v_474_0;
  wire [2:0] v_475_0;
  wire [0:0] v_476_0;
  wire [2:0] v_477_0;
  wire [2:0] v_478_0;
  wire [2:0] v_479_0;
  wire [2:0] v_480_0;
  wire [2:0] v_481_0;
  wire [2:0] v_482_0;
  wire [2:0] v_483_0;
  wire [2:0] v_484_0;
  wire [2:0] v_485_0;
  wire [2:0] v_486_0;
  wire [2:0] v_487_0;
  wire [2:0] v_488_0;
  wire [2:0] v_489_0;
  wire [0:0] v_490_0;
  wire [2:0] v_491_0;
  wire [2:0] v_491_1;
  wire [4:0] v_492_0;
  wire [4:0] v_493_0;
  wire [4:0] v_494_0;
  wire [0:0] v_495_0;
  wire [2:0] v_496_0;
  wire [0:0] v_497_0;
  wire [0:0] v_498_0;
  wire [0:0] v_499_0;
  wire [4:0] v_500_0;
  wire [4:0] v_501_0;
  wire [4:0] v_502_0;
  wire [0:0] v_503_0;
  wire [2:0] v_504_0;
  wire [2:0] v_505_0;
  wire [2:0] v_506_0;
  wire [0:0] v_507_0;
  wire [0:0] v_508_0;
  wire [0:0] v_509_0;
  wire [0:0] v_510_0;
  wire [0:0] v_511_0;
  wire [2:0] v_512_0;
  wire [0:0] v_513_0;
  reg [2:0] v_514_0 = 3'h0;
  wire [0:0] v_515_0;
  wire [0:0] v_516_0;
  wire [0:0] v_517_0;
  wire [0:0] v_518_0;
  wire [0:0] v_519_0;
  wire [0:0] v_520_0;
  wire [0:0] v_521_0;
  wire [0:0] v_522_0;
  wire [0:0] v_523_0;
  wire [0:0] v_524_0;
  wire [0:0] v_525_0;
  wire [0:0] v_526_0;
  wire [0:0] v_527_0;
  wire [0:0] v_528_0;
  wire [0:0] v_529_0;
  wire [0:0] v_530_0;
  wire [0:0] v_531_0;
  wire [0:0] v_532_0;
  wire [0:0] v_533_0;
  wire [0:0] v_534_0;
  wire [0:0] v_535_0;
  wire [0:0] v_536_0;
  wire [0:0] v_537_0;
  wire [0:0] v_538_0;
  wire [0:0] v_539_0;
  wire [0:0] v_540_0;
  wire [0:0] v_541_0;
  wire [0:0] v_542_0;
  wire [0:0] v_543_0;
  wire [2:0] v_544_0;
  wire [2:0] v_545_0;
  wire [2:0] v_546_0;
  wire [2:0] v_547_0;
  wire [2:0] v_548_0;
  wire [2:0] v_549_0;
  wire [2:0] v_550_0;
  wire [2:0] v_551_0;
  wire [2:0] v_552_0;
  wire [2:0] v_553_0;
  wire [2:0] v_554_0;
  wire [2:0] v_555_0;
  wire [2:0] v_556_0;
  wire [2:0] v_557_0;
  wire [2:0] v_558_0;
  wire [2:0] v_559_0;
  wire [2:0] v_560_0;
  wire [2:0] v_561_0;
  wire [2:0] v_562_0;
  wire [0:0] v_563_0;
  wire [0:0] v_564_0;
  wire [15:0] v_565_0;
  wire [0:0] v_566_0;
  wire [0:0] v_567_0;
  wire [0:0] v_568_0;
  wire [0:0] v_569_0;
  wire [0:0] v_570_0;
  wire [0:0] v_571_0;
  wire [0:0] v_572_0;
  wire [0:0] v_573_0;
  wire [0:0] v_574_0;
  wire [0:0] v_575_0;
  wire [0:0] v_576_0;
  wire [0:0] v_577_0;
  reg [15:0] v_578_0 = 16'h0;
  wire [0:0] v_579_0;
  wire [0:0] v_580_0;
  wire [0:0] v_581_0;
  wire [0:0] v_582_0;
  wire [0:0] v_583_0;
  wire [0:0] v_584_0;
  wire [0:0] v_585_0;
  wire [0:0] v_586_0;
  wire [0:0] v_587_0;
  wire [0:0] v_588_0;
  wire [0:0] v_589_0;
  wire [0:0] v_590_0;
  wire [0:0] v_591_0;
  wire [0:0] v_592_0;
  wire [0:0] v_593_0;
  wire [0:0] v_594_0;
  wire [0:0] v_595_0;
  wire [0:0] v_596_0;
  reg [9:0] v_597_0 = 10'h0;
  wire [0:0] v_598_0;
  wire [0:0] v_599_0;
  wire [0:0] v_600_0;
  wire [0:0] v_601_0;
  wire [0:0] v_602_0;
  wire [0:0] v_603_0;
  wire [0:0] v_604_0;
  wire [0:0] v_605_0;
  wire [0:0] v_606_0;
  wire [0:0] v_607_0;
  wire [0:0] v_608_0;
  wire [0:0] v_609_0;
  wire [0:0] v_610_0;
  wire [0:0] v_611_0;
  wire [0:0] v_612_0;
  wire [0:0] v_613_0;
  wire [0:0] v_614_0;
  reg [0:0] v_615_0 = 1'h0;
  reg [0:0] v_616_0 = 1'h0;
  wire [0:0] v_617_0;
  wire [0:0] v_618_0;
  wire [0:0] v_619_0;
  reg [0:0] v_620_0 = 1'h0;
  wire [0:0] v_621_0;
  wire [0:0] v_622_0;
  wire [0:0] v_623_0;
  wire [0:0] v_624_0;
  wire [0:0] v_625_0;
  wire [0:0] v_626_0;
  wire [0:0] v_627_0;
  wire [0:0] v_628_0;
  wire [0:0] v_629_0;
  wire [0:0] v_630_0;
  wire [0:0] v_631_0;
  wire [0:0] v_632_0;
  wire [0:0] v_633_0;
  wire [0:0] v_634_0;
  wire [0:0] v_635_0;
  wire [0:0] v_636_0;
  wire [0:0] v_637_0;
  wire [0:0] v_638_0;
  wire [0:0] v_639_0;
  wire [0:0] v_640_0;
  wire [0:0] v_641_0;
  reg [0:0] v_642_0 = 1'h0;
  wire [0:0] v_643_0;
  wire [0:0] v_644_0;
  wire [0:0] v_645_0;
  wire [0:0] v_646_0;
  wire [0:0] v_647_0;
  wire [0:0] v_648_0;
  wire [0:0] v_649_0;
  wire [0:0] v_650_0;
  wire [0:0] v_651_0;
  wire [0:0] v_652_0;
  wire [0:0] v_653_0;
  wire [0:0] v_654_0;
  wire [0:0] v_655_0;
  wire [0:0] v_656_0;
  wire [9:0] v_657_0;
  wire [9:0] v_658_0;
  wire [9:0] v_659_0;
  wire [9:0] v_660_0;
  wire [9:0] v_661_0;
  wire [9:0] v_662_0;
  wire [9:0] v_663_0;
  wire [9:0] v_664_0;
  wire [9:0] v_665_0;
  wire [9:0] v_666_0;
  wire [9:0] v_667_0;
  wire [9:0] v_668_0;
  wire [9:0] v_669_0;
  wire [9:0] v_670_0;
  wire [9:0] v_671_0;
  wire [9:0] v_672_0;
  wire [9:0] v_673_0;
  wire [9:0] v_674_0;
  wire [0:0] v_675_0;
  wire [9:0] v_676_0;
  wire [9:0] v_677_0;
  wire [9:0] v_678_0;
  wire [9:0] v_679_0;
  wire [9:0] v_680_0;
  wire [9:0] v_681_0;
  wire [9:0] v_682_0;
  wire [9:0] v_683_0;
  wire [9:0] v_684_0;
  wire [9:0] v_685_0;
  wire [9:0] v_686_0;
  wire [9:0] v_687_0;
  wire [9:0] v_688_0;
  wire [0:0] v_689_0;
  reg [2:0] v_690_0 = 3'h0;
  wire [0:0] v_691_0;
  wire [0:0] v_692_0;
  wire [0:0] v_693_0;
  wire [2:0] v_694_0;
  wire [2:0] v_695_0;
  wire [2:0] v_696_0;
  reg [2:0] v_697_0 = 3'h0;
  wire [0:0] v_698_0;
  wire [0:0] v_699_0;
  wire [0:0] v_700_0;
  wire [2:0] v_701_0;
  wire [2:0] v_702_0;
  wire [2:0] v_703_0;
  reg [2:0] v_704_0 = 3'h0;
  wire [0:0] v_705_0;
  wire [0:0] v_706_0;
  wire [0:0] v_707_0;
  wire [2:0] v_708_0;
  wire [2:0] v_709_0;
  wire [2:0] v_710_0;
  reg [2:0] v_711_0 = 3'h0;
  wire [0:0] v_712_0;
  wire [0:0] v_713_0;
  wire [0:0] v_714_0;
  wire [2:0] v_715_0;
  wire [2:0] v_716_0;
  wire [2:0] v_717_0;
  reg [2:0] v_718_0 = 3'h0;
  wire [0:0] v_719_0;
  wire [0:0] v_720_0;
  wire [0:0] v_721_0;
  wire [2:0] v_722_0;
  wire [2:0] v_723_0;
  wire [2:0] v_724_0;
  reg [2:0] v_725_0 = 3'h0;
  wire [0:0] v_726_0;
  wire [0:0] v_727_0;
  wire [0:0] v_728_0;
  wire [2:0] v_729_0;
  wire [2:0] v_730_0;
  wire [2:0] v_731_0;
  reg [2:0] v_732_0 = 3'h0;
  wire [0:0] v_733_0;
  wire [0:0] v_734_0;
  wire [0:0] v_735_0;
  wire [2:0] v_736_0;
  wire [2:0] v_737_0;
  wire [2:0] v_738_0;
  reg [2:0] v_739_0 = 3'h0;
  wire [0:0] v_740_0;
  wire [0:0] v_741_0;
  wire [0:0] v_742_0;
  wire [2:0] v_743_0;
  wire [2:0] v_744_0;
  wire [2:0] v_745_0;
  reg [2:0] v_746_0 = 3'h0;
  wire [0:0] v_747_0;
  wire [0:0] v_748_0;
  wire [0:0] v_749_0;
  wire [2:0] v_750_0;
  wire [2:0] v_751_0;
  wire [2:0] v_752_0;
  reg [2:0] v_753_0 = 3'h0;
  wire [0:0] v_754_0;
  wire [0:0] v_755_0;
  wire [0:0] v_756_0;
  wire [2:0] v_757_0;
  wire [2:0] v_758_0;
  wire [2:0] v_759_0;
  reg [2:0] v_760_0 = 3'h0;
  wire [0:0] v_761_0;
  wire [0:0] v_762_0;
  wire [0:0] v_763_0;
  wire [2:0] v_764_0;
  wire [2:0] v_765_0;
  wire [2:0] v_766_0;
  reg [2:0] v_767_0 = 3'h0;
  wire [0:0] v_768_0;
  wire [0:0] v_769_0;
  wire [0:0] v_770_0;
  wire [2:0] v_771_0;
  wire [2:0] v_772_0;
  wire [2:0] v_773_0;
  reg [2:0] v_774_0 = 3'h0;
  wire [0:0] v_775_0;
  wire [0:0] v_776_0;
  wire [0:0] v_777_0;
  wire [2:0] v_778_0;
  wire [2:0] v_779_0;
  wire [2:0] v_780_0;
  reg [2:0] v_781_0 = 3'h0;
  wire [0:0] v_782_0;
  wire [0:0] v_783_0;
  wire [0:0] v_784_0;
  wire [2:0] v_785_0;
  wire [2:0] v_786_0;
  wire [2:0] v_787_0;
  reg [2:0] v_788_0 = 3'h0;
  wire [0:0] v_789_0;
  wire [0:0] v_790_0;
  wire [0:0] v_791_0;
  wire [2:0] v_792_0;
  wire [2:0] v_793_0;
  wire [2:0] v_794_0;
  reg [2:0] v_795_0 = 3'h0;
  wire [0:0] v_796_0;
  wire [0:0] v_797_0;
  wire [0:0] v_798_0;
  wire [2:0] v_799_0;
  wire [2:0] v_800_0;
  wire [2:0] v_801_0;
  reg [2:0] v_802_0 = 3'h0;
  wire [0:0] v_803_0;
  wire [0:0] v_804_0;
  wire [0:0] v_805_0;
  wire [2:0] v_806_0;
  wire [2:0] v_807_0;
  wire [2:0] v_808_0;
  reg [2:0] v_809_0 = 3'h0;
  wire [0:0] v_810_0;
  wire [0:0] v_811_0;
  wire [0:0] v_812_0;
  wire [2:0] v_813_0;
  wire [2:0] v_814_0;
  wire [2:0] v_815_0;
  reg [2:0] v_816_0 = 3'h0;
  wire [0:0] v_817_0;
  wire [0:0] v_818_0;
  wire [0:0] v_819_0;
  wire [2:0] v_820_0;
  wire [2:0] v_821_0;
  wire [2:0] v_822_0;
  reg [2:0] v_823_0 = 3'h0;
  wire [0:0] v_824_0;
  wire [0:0] v_825_0;
  wire [0:0] v_826_0;
  wire [2:0] v_827_0;
  wire [2:0] v_828_0;
  wire [2:0] v_829_0;
  reg [2:0] v_830_0 = 3'h0;
  wire [0:0] v_831_0;
  wire [0:0] v_832_0;
  wire [0:0] v_833_0;
  wire [2:0] v_834_0;
  wire [2:0] v_835_0;
  wire [2:0] v_836_0;
  reg [2:0] v_837_0 = 3'h0;
  wire [0:0] v_838_0;
  wire [0:0] v_839_0;
  wire [0:0] v_840_0;
  wire [2:0] v_841_0;
  wire [2:0] v_842_0;
  wire [2:0] v_843_0;
  reg [2:0] v_844_0 = 3'h0;
  wire [0:0] v_845_0;
  wire [0:0] v_846_0;
  wire [0:0] v_847_0;
  wire [2:0] v_848_0;
  wire [2:0] v_849_0;
  wire [2:0] v_850_0;
  reg [2:0] v_851_0 = 3'h0;
  wire [0:0] v_852_0;
  wire [0:0] v_853_0;
  wire [0:0] v_854_0;
  wire [2:0] v_855_0;
  wire [2:0] v_856_0;
  wire [2:0] v_857_0;
  reg [2:0] v_858_0 = 3'h0;
  wire [0:0] v_859_0;
  wire [0:0] v_860_0;
  wire [0:0] v_861_0;
  wire [2:0] v_862_0;
  wire [2:0] v_863_0;
  wire [2:0] v_864_0;
  reg [2:0] v_865_0 = 3'h0;
  wire [0:0] v_866_0;
  wire [0:0] v_867_0;
  wire [0:0] v_868_0;
  wire [2:0] v_869_0;
  wire [2:0] v_870_0;
  wire [2:0] v_871_0;
  reg [2:0] v_872_0 = 3'h0;
  wire [0:0] v_873_0;
  wire [0:0] v_874_0;
  wire [0:0] v_875_0;
  wire [2:0] v_876_0;
  wire [2:0] v_877_0;
  wire [2:0] v_878_0;
  reg [2:0] v_879_0 = 3'h0;
  wire [0:0] v_880_0;
  wire [0:0] v_881_0;
  wire [0:0] v_882_0;
  wire [2:0] v_883_0;
  wire [2:0] v_884_0;
  wire [2:0] v_885_0;
  reg [2:0] v_886_0 = 3'h0;
  wire [0:0] v_887_0;
  wire [0:0] v_888_0;
  wire [0:0] v_889_0;
  wire [2:0] v_890_0;
  wire [2:0] v_891_0;
  wire [2:0] v_892_0;
  reg [2:0] v_893_0 = 3'h0;
  wire [0:0] v_894_0;
  wire [0:0] v_895_0;
  wire [0:0] v_896_0;
  wire [2:0] v_897_0;
  wire [2:0] v_898_0;
  wire [2:0] v_899_0;
  reg [2:0] v_900_0 = 3'h0;
  wire [0:0] v_901_0;
  wire [0:0] v_902_0;
  wire [0:0] v_903_0;
  wire [2:0] v_904_0;
  wire [2:0] v_905_0;
  wire [2:0] v_906_0;
  reg [2:0] v_907_0 = 3'h0;
  wire [0:0] v_908_0;
  wire [0:0] v_909_0;
  wire [0:0] v_910_0;
  wire [2:0] v_911_0;
  wire [2:0] v_912_0;
  wire [2:0] v_913_0;
  reg [2:0] v_914_0 = 3'h0;
  wire [0:0] v_915_0;
  wire [0:0] v_916_0;
  wire [0:0] v_917_0;
  wire [2:0] v_918_0;
  wire [2:0] v_919_0;
  wire [2:0] v_920_0;
  reg [2:0] v_921_0 = 3'h0;
  wire [0:0] v_922_0;
  wire [0:0] v_923_0;
  wire [0:0] v_924_0;
  wire [2:0] v_925_0;
  wire [2:0] v_926_0;
  wire [2:0] v_927_0;
  reg [2:0] v_928_0 = 3'h0;
  wire [0:0] v_929_0;
  wire [0:0] v_930_0;
  wire [0:0] v_931_0;
  wire [2:0] v_932_0;
  wire [2:0] v_933_0;
  wire [2:0] v_934_0;
  reg [2:0] v_935_0 = 3'h0;
  wire [0:0] v_936_0;
  wire [0:0] v_937_0;
  wire [0:0] v_938_0;
  wire [2:0] v_939_0;
  wire [2:0] v_940_0;
  wire [2:0] v_941_0;
  reg [2:0] v_942_0 = 3'h0;
  wire [0:0] v_943_0;
  wire [0:0] v_944_0;
  wire [0:0] v_945_0;
  wire [2:0] v_946_0;
  wire [2:0] v_947_0;
  wire [2:0] v_948_0;
  reg [2:0] v_949_0 = 3'h0;
  wire [0:0] v_950_0;
  wire [0:0] v_951_0;
  wire [0:0] v_952_0;
  wire [2:0] v_953_0;
  wire [2:0] v_954_0;
  wire [2:0] v_955_0;
  reg [2:0] v_956_0 = 3'h0;
  wire [0:0] v_957_0;
  wire [0:0] v_958_0;
  wire [0:0] v_959_0;
  wire [2:0] v_960_0;
  wire [2:0] v_961_0;
  wire [2:0] v_962_0;
  reg [2:0] v_963_0 = 3'h0;
  wire [0:0] v_964_0;
  wire [0:0] v_965_0;
  wire [0:0] v_966_0;
  wire [2:0] v_967_0;
  wire [2:0] v_968_0;
  wire [2:0] v_969_0;
  reg [2:0] v_970_0 = 3'h0;
  wire [0:0] v_971_0;
  wire [0:0] v_972_0;
  wire [0:0] v_973_0;
  wire [2:0] v_974_0;
  wire [2:0] v_975_0;
  wire [2:0] v_976_0;
  reg [2:0] v_977_0 = 3'h0;
  wire [0:0] v_978_0;
  wire [0:0] v_979_0;
  wire [0:0] v_980_0;
  wire [2:0] v_981_0;
  wire [2:0] v_982_0;
  wire [2:0] v_983_0;
  reg [2:0] v_984_0 = 3'h0;
  wire [0:0] v_985_0;
  wire [0:0] v_986_0;
  wire [0:0] v_987_0;
  wire [2:0] v_988_0;
  wire [2:0] v_989_0;
  wire [2:0] v_990_0;
  reg [2:0] v_991_0 = 3'h0;
  wire [0:0] v_992_0;
  wire [0:0] v_993_0;
  wire [0:0] v_994_0;
  wire [2:0] v_995_0;
  wire [2:0] v_996_0;
  wire [2:0] v_997_0;
  reg [2:0] v_998_0 = 3'h0;
  wire [0:0] v_999_0;
  wire [0:0] v_1000_0;
  wire [0:0] v_1001_0;
  wire [2:0] v_1002_0;
  wire [2:0] v_1003_0;
  wire [2:0] v_1004_0;
  reg [2:0] v_1005_0 = 3'h0;
  wire [0:0] v_1006_0;
  wire [0:0] v_1007_0;
  wire [0:0] v_1008_0;
  wire [2:0] v_1009_0;
  wire [2:0] v_1010_0;
  wire [2:0] v_1011_0;
  reg [2:0] v_1012_0 = 3'h0;
  wire [0:0] v_1013_0;
  wire [0:0] v_1014_0;
  wire [0:0] v_1015_0;
  wire [2:0] v_1016_0;
  wire [2:0] v_1017_0;
  wire [2:0] v_1018_0;
  reg [2:0] v_1019_0 = 3'h0;
  wire [0:0] v_1020_0;
  wire [0:0] v_1021_0;
  wire [0:0] v_1022_0;
  wire [2:0] v_1023_0;
  wire [2:0] v_1024_0;
  wire [2:0] v_1025_0;
  reg [2:0] v_1026_0 = 3'h0;
  wire [0:0] v_1027_0;
  wire [0:0] v_1028_0;
  wire [0:0] v_1029_0;
  wire [2:0] v_1030_0;
  wire [2:0] v_1031_0;
  wire [2:0] v_1032_0;
  reg [2:0] v_1033_0 = 3'h0;
  wire [0:0] v_1034_0;
  wire [0:0] v_1035_0;
  wire [0:0] v_1036_0;
  wire [2:0] v_1037_0;
  wire [2:0] v_1038_0;
  wire [2:0] v_1039_0;
  reg [2:0] v_1040_0 = 3'h0;
  wire [0:0] v_1041_0;
  wire [0:0] v_1042_0;
  wire [0:0] v_1043_0;
  wire [2:0] v_1044_0;
  wire [2:0] v_1045_0;
  wire [2:0] v_1046_0;
  reg [2:0] v_1047_0 = 3'h0;
  wire [0:0] v_1048_0;
  wire [0:0] v_1049_0;
  wire [0:0] v_1050_0;
  wire [2:0] v_1051_0;
  wire [2:0] v_1052_0;
  wire [2:0] v_1053_0;
  reg [2:0] v_1054_0 = 3'h0;
  wire [0:0] v_1055_0;
  wire [0:0] v_1056_0;
  wire [0:0] v_1057_0;
  wire [2:0] v_1058_0;
  wire [2:0] v_1059_0;
  wire [2:0] v_1060_0;
  reg [2:0] v_1061_0 = 3'h0;
  wire [0:0] v_1062_0;
  wire [0:0] v_1063_0;
  wire [0:0] v_1064_0;
  wire [2:0] v_1065_0;
  wire [2:0] v_1066_0;
  wire [2:0] v_1067_0;
  reg [2:0] v_1068_0 = 3'h0;
  wire [0:0] v_1069_0;
  wire [0:0] v_1070_0;
  wire [0:0] v_1071_0;
  wire [2:0] v_1072_0;
  wire [2:0] v_1073_0;
  wire [2:0] v_1074_0;
  reg [2:0] v_1075_0 = 3'h0;
  wire [0:0] v_1076_0;
  wire [0:0] v_1077_0;
  wire [0:0] v_1078_0;
  wire [2:0] v_1079_0;
  wire [2:0] v_1080_0;
  wire [2:0] v_1081_0;
  reg [2:0] v_1082_0 = 3'h0;
  wire [0:0] v_1083_0;
  wire [0:0] v_1084_0;
  wire [0:0] v_1085_0;
  wire [2:0] v_1086_0;
  wire [2:0] v_1087_0;
  wire [2:0] v_1088_0;
  reg [2:0] v_1089_0 = 3'h0;
  wire [0:0] v_1090_0;
  wire [0:0] v_1091_0;
  wire [0:0] v_1092_0;
  wire [2:0] v_1093_0;
  wire [2:0] v_1094_0;
  wire [2:0] v_1095_0;
  reg [2:0] v_1096_0 = 3'h0;
  wire [0:0] v_1097_0;
  wire [0:0] v_1098_0;
  wire [0:0] v_1099_0;
  wire [2:0] v_1100_0;
  wire [2:0] v_1101_0;
  wire [2:0] v_1102_0;
  reg [2:0] v_1103_0 = 3'h0;
  wire [0:0] v_1104_0;
  wire [0:0] v_1105_0;
  wire [0:0] v_1106_0;
  wire [2:0] v_1107_0;
  wire [2:0] v_1108_0;
  wire [2:0] v_1109_0;
  reg [2:0] v_1110_0 = 3'h0;
  wire [0:0] v_1111_0;
  wire [0:0] v_1112_0;
  wire [0:0] v_1113_0;
  wire [2:0] v_1114_0;
  wire [2:0] v_1115_0;
  wire [2:0] v_1116_0;
  reg [2:0] v_1117_0 = 3'h0;
  wire [0:0] v_1118_0;
  wire [0:0] v_1119_0;
  wire [0:0] v_1120_0;
  wire [2:0] v_1121_0;
  wire [2:0] v_1122_0;
  wire [2:0] v_1123_0;
  reg [2:0] v_1124_0 = 3'h0;
  wire [0:0] v_1125_0;
  wire [0:0] v_1126_0;
  wire [0:0] v_1127_0;
  wire [2:0] v_1128_0;
  wire [2:0] v_1129_0;
  wire [2:0] v_1130_0;
  reg [2:0] v_1131_0 = 3'h0;
  wire [0:0] v_1132_0;
  wire [0:0] v_1133_0;
  wire [0:0] v_1134_0;
  wire [2:0] v_1135_0;
  wire [2:0] v_1136_0;
  wire [2:0] v_1137_0;
  reg [2:0] v_1138_0 = 3'h0;
  wire [0:0] v_1139_0;
  wire [0:0] v_1140_0;
  wire [0:0] v_1141_0;
  wire [2:0] v_1142_0;
  wire [2:0] v_1143_0;
  wire [2:0] v_1144_0;
  reg [2:0] v_1145_0 = 3'h0;
  wire [0:0] v_1146_0;
  wire [0:0] v_1147_0;
  wire [0:0] v_1148_0;
  wire [2:0] v_1149_0;
  wire [2:0] v_1150_0;
  wire [2:0] v_1151_0;
  reg [2:0] v_1152_0 = 3'h0;
  wire [0:0] v_1153_0;
  wire [0:0] v_1154_0;
  wire [0:0] v_1155_0;
  wire [2:0] v_1156_0;
  wire [2:0] v_1157_0;
  wire [2:0] v_1158_0;
  reg [2:0] v_1159_0 = 3'h0;
  wire [0:0] v_1160_0;
  wire [0:0] v_1161_0;
  wire [0:0] v_1162_0;
  wire [2:0] v_1163_0;
  wire [2:0] v_1164_0;
  wire [2:0] v_1165_0;
  reg [2:0] v_1166_0 = 3'h0;
  wire [0:0] v_1167_0;
  wire [0:0] v_1168_0;
  wire [0:0] v_1169_0;
  wire [2:0] v_1170_0;
  wire [2:0] v_1171_0;
  wire [2:0] v_1172_0;
  reg [2:0] v_1173_0 = 3'h0;
  wire [0:0] v_1174_0;
  wire [0:0] v_1175_0;
  wire [0:0] v_1176_0;
  wire [2:0] v_1177_0;
  wire [2:0] v_1178_0;
  wire [2:0] v_1179_0;
  reg [2:0] v_1180_0 = 3'h0;
  wire [0:0] v_1181_0;
  wire [0:0] v_1182_0;
  wire [0:0] v_1183_0;
  wire [2:0] v_1184_0;
  wire [2:0] v_1185_0;
  wire [2:0] v_1186_0;
  reg [2:0] v_1187_0 = 3'h0;
  wire [0:0] v_1188_0;
  wire [0:0] v_1189_0;
  wire [0:0] v_1190_0;
  wire [2:0] v_1191_0;
  wire [2:0] v_1192_0;
  wire [2:0] v_1193_0;
  reg [2:0] v_1194_0 = 3'h0;
  wire [0:0] v_1195_0;
  wire [0:0] v_1196_0;
  wire [0:0] v_1197_0;
  wire [2:0] v_1198_0;
  wire [2:0] v_1199_0;
  wire [2:0] v_1200_0;
  reg [2:0] v_1201_0 = 3'h0;
  wire [0:0] v_1202_0;
  wire [0:0] v_1203_0;
  wire [0:0] v_1204_0;
  wire [2:0] v_1205_0;
  wire [2:0] v_1206_0;
  wire [2:0] v_1207_0;
  reg [2:0] v_1208_0 = 3'h0;
  wire [0:0] v_1209_0;
  wire [0:0] v_1210_0;
  wire [0:0] v_1211_0;
  wire [2:0] v_1212_0;
  wire [2:0] v_1213_0;
  wire [2:0] v_1214_0;
  reg [2:0] v_1215_0 = 3'h0;
  wire [0:0] v_1216_0;
  wire [0:0] v_1217_0;
  wire [0:0] v_1218_0;
  wire [2:0] v_1219_0;
  wire [2:0] v_1220_0;
  wire [2:0] v_1221_0;
  reg [2:0] v_1222_0 = 3'h0;
  wire [0:0] v_1223_0;
  wire [0:0] v_1224_0;
  wire [0:0] v_1225_0;
  wire [2:0] v_1226_0;
  wire [2:0] v_1227_0;
  wire [2:0] v_1228_0;
  reg [2:0] v_1229_0 = 3'h0;
  wire [0:0] v_1230_0;
  wire [0:0] v_1231_0;
  wire [0:0] v_1232_0;
  wire [2:0] v_1233_0;
  wire [2:0] v_1234_0;
  wire [2:0] v_1235_0;
  reg [2:0] v_1236_0 = 3'h0;
  wire [0:0] v_1237_0;
  wire [0:0] v_1238_0;
  wire [0:0] v_1239_0;
  wire [2:0] v_1240_0;
  wire [2:0] v_1241_0;
  wire [2:0] v_1242_0;
  reg [2:0] v_1243_0 = 3'h0;
  wire [0:0] v_1244_0;
  wire [0:0] v_1245_0;
  wire [0:0] v_1246_0;
  wire [2:0] v_1247_0;
  wire [2:0] v_1248_0;
  wire [2:0] v_1249_0;
  reg [2:0] v_1250_0 = 3'h0;
  wire [0:0] v_1251_0;
  wire [0:0] v_1252_0;
  wire [0:0] v_1253_0;
  wire [2:0] v_1254_0;
  wire [2:0] v_1255_0;
  wire [2:0] v_1256_0;
  reg [2:0] v_1257_0 = 3'h0;
  wire [0:0] v_1258_0;
  wire [0:0] v_1259_0;
  wire [0:0] v_1260_0;
  wire [2:0] v_1261_0;
  wire [2:0] v_1262_0;
  wire [2:0] v_1263_0;
  reg [2:0] v_1264_0 = 3'h0;
  wire [0:0] v_1265_0;
  wire [0:0] v_1266_0;
  wire [0:0] v_1267_0;
  wire [2:0] v_1268_0;
  wire [2:0] v_1269_0;
  wire [2:0] v_1270_0;
  reg [2:0] v_1271_0 = 3'h0;
  wire [0:0] v_1272_0;
  wire [0:0] v_1273_0;
  wire [0:0] v_1274_0;
  wire [2:0] v_1275_0;
  wire [2:0] v_1276_0;
  wire [2:0] v_1277_0;
  reg [2:0] v_1278_0 = 3'h0;
  wire [0:0] v_1279_0;
  wire [0:0] v_1280_0;
  wire [0:0] v_1281_0;
  wire [2:0] v_1282_0;
  wire [2:0] v_1283_0;
  wire [2:0] v_1284_0;
  reg [2:0] v_1285_0 = 3'h0;
  wire [0:0] v_1286_0;
  wire [0:0] v_1287_0;
  wire [0:0] v_1288_0;
  wire [2:0] v_1289_0;
  wire [2:0] v_1290_0;
  wire [2:0] v_1291_0;
  reg [2:0] v_1292_0 = 3'h0;
  wire [0:0] v_1293_0;
  wire [0:0] v_1294_0;
  wire [0:0] v_1295_0;
  wire [2:0] v_1296_0;
  wire [2:0] v_1297_0;
  wire [2:0] v_1298_0;
  reg [2:0] v_1299_0 = 3'h0;
  wire [0:0] v_1300_0;
  wire [0:0] v_1301_0;
  wire [0:0] v_1302_0;
  wire [2:0] v_1303_0;
  wire [2:0] v_1304_0;
  wire [2:0] v_1305_0;
  reg [2:0] v_1306_0 = 3'h0;
  wire [0:0] v_1307_0;
  wire [0:0] v_1308_0;
  wire [0:0] v_1309_0;
  wire [2:0] v_1310_0;
  wire [2:0] v_1311_0;
  wire [2:0] v_1312_0;
  reg [2:0] v_1313_0 = 3'h0;
  wire [0:0] v_1314_0;
  wire [0:0] v_1315_0;
  wire [0:0] v_1316_0;
  wire [2:0] v_1317_0;
  wire [2:0] v_1318_0;
  wire [2:0] v_1319_0;
  reg [2:0] v_1320_0 = 3'h0;
  wire [0:0] v_1321_0;
  wire [0:0] v_1322_0;
  wire [0:0] v_1323_0;
  wire [2:0] v_1324_0;
  wire [2:0] v_1325_0;
  wire [2:0] v_1326_0;
  reg [2:0] v_1327_0 = 3'h0;
  wire [0:0] v_1328_0;
  wire [0:0] v_1329_0;
  wire [0:0] v_1330_0;
  wire [2:0] v_1331_0;
  wire [2:0] v_1332_0;
  wire [2:0] v_1333_0;
  reg [2:0] v_1334_0 = 3'h0;
  wire [0:0] v_1335_0;
  wire [0:0] v_1336_0;
  wire [0:0] v_1337_0;
  wire [2:0] v_1338_0;
  wire [2:0] v_1339_0;
  wire [2:0] v_1340_0;
  reg [2:0] v_1341_0 = 3'h0;
  wire [0:0] v_1342_0;
  wire [0:0] v_1343_0;
  wire [0:0] v_1344_0;
  wire [2:0] v_1345_0;
  wire [2:0] v_1346_0;
  wire [2:0] v_1347_0;
  reg [2:0] v_1348_0 = 3'h0;
  wire [0:0] v_1349_0;
  wire [0:0] v_1350_0;
  wire [0:0] v_1351_0;
  wire [2:0] v_1352_0;
  wire [2:0] v_1353_0;
  wire [2:0] v_1354_0;
  reg [2:0] v_1355_0 = 3'h0;
  wire [0:0] v_1356_0;
  wire [0:0] v_1357_0;
  wire [0:0] v_1358_0;
  wire [2:0] v_1359_0;
  wire [2:0] v_1360_0;
  wire [2:0] v_1361_0;
  reg [2:0] v_1362_0 = 3'h0;
  wire [0:0] v_1363_0;
  wire [0:0] v_1364_0;
  wire [0:0] v_1365_0;
  wire [2:0] v_1366_0;
  wire [2:0] v_1367_0;
  wire [2:0] v_1368_0;
  reg [2:0] v_1369_0 = 3'h0;
  wire [0:0] v_1370_0;
  wire [0:0] v_1371_0;
  wire [0:0] v_1372_0;
  wire [2:0] v_1373_0;
  wire [2:0] v_1374_0;
  wire [2:0] v_1375_0;
  reg [2:0] v_1376_0 = 3'h0;
  wire [0:0] v_1377_0;
  wire [0:0] v_1378_0;
  wire [0:0] v_1379_0;
  wire [2:0] v_1380_0;
  wire [2:0] v_1381_0;
  wire [2:0] v_1382_0;
  reg [2:0] v_1383_0 = 3'h0;
  wire [0:0] v_1384_0;
  wire [0:0] v_1385_0;
  wire [0:0] v_1386_0;
  wire [2:0] v_1387_0;
  wire [2:0] v_1388_0;
  wire [2:0] v_1389_0;
  reg [2:0] v_1390_0 = 3'h0;
  wire [0:0] v_1391_0;
  wire [0:0] v_1392_0;
  wire [0:0] v_1393_0;
  wire [2:0] v_1394_0;
  wire [2:0] v_1395_0;
  wire [2:0] v_1396_0;
  reg [2:0] v_1397_0 = 3'h0;
  wire [0:0] v_1398_0;
  wire [0:0] v_1399_0;
  wire [0:0] v_1400_0;
  wire [2:0] v_1401_0;
  wire [2:0] v_1402_0;
  wire [2:0] v_1403_0;
  reg [2:0] v_1404_0 = 3'h0;
  wire [0:0] v_1405_0;
  wire [0:0] v_1406_0;
  wire [0:0] v_1407_0;
  wire [2:0] v_1408_0;
  wire [2:0] v_1409_0;
  wire [2:0] v_1410_0;
  reg [2:0] v_1411_0 = 3'h0;
  wire [0:0] v_1412_0;
  wire [0:0] v_1413_0;
  wire [0:0] v_1414_0;
  wire [2:0] v_1415_0;
  wire [2:0] v_1416_0;
  wire [2:0] v_1417_0;
  reg [2:0] v_1418_0 = 3'h0;
  wire [0:0] v_1419_0;
  wire [0:0] v_1420_0;
  wire [0:0] v_1421_0;
  wire [2:0] v_1422_0;
  wire [2:0] v_1423_0;
  wire [2:0] v_1424_0;
  reg [2:0] v_1425_0 = 3'h0;
  wire [0:0] v_1426_0;
  wire [0:0] v_1427_0;
  wire [0:0] v_1428_0;
  wire [2:0] v_1429_0;
  wire [2:0] v_1430_0;
  wire [2:0] v_1431_0;
  reg [2:0] v_1432_0 = 3'h0;
  wire [0:0] v_1433_0;
  wire [0:0] v_1434_0;
  wire [0:0] v_1435_0;
  wire [2:0] v_1436_0;
  wire [2:0] v_1437_0;
  wire [2:0] v_1438_0;
  reg [2:0] v_1439_0 = 3'h0;
  wire [0:0] v_1440_0;
  wire [0:0] v_1441_0;
  wire [0:0] v_1442_0;
  wire [2:0] v_1443_0;
  wire [2:0] v_1444_0;
  wire [2:0] v_1445_0;
  reg [2:0] v_1446_0 = 3'h0;
  wire [0:0] v_1447_0;
  wire [0:0] v_1448_0;
  wire [0:0] v_1449_0;
  wire [2:0] v_1450_0;
  wire [2:0] v_1451_0;
  wire [2:0] v_1452_0;
  reg [2:0] v_1453_0 = 3'h0;
  wire [0:0] v_1454_0;
  wire [0:0] v_1455_0;
  wire [0:0] v_1456_0;
  wire [2:0] v_1457_0;
  wire [2:0] v_1458_0;
  wire [2:0] v_1459_0;
  reg [2:0] v_1460_0 = 3'h0;
  wire [0:0] v_1461_0;
  wire [0:0] v_1462_0;
  wire [0:0] v_1463_0;
  wire [2:0] v_1464_0;
  wire [2:0] v_1465_0;
  wire [2:0] v_1466_0;
  reg [2:0] v_1467_0 = 3'h0;
  wire [0:0] v_1468_0;
  wire [0:0] v_1469_0;
  wire [0:0] v_1470_0;
  wire [2:0] v_1471_0;
  wire [2:0] v_1472_0;
  wire [2:0] v_1473_0;
  reg [2:0] v_1474_0 = 3'h0;
  wire [0:0] v_1475_0;
  wire [0:0] v_1476_0;
  wire [0:0] v_1477_0;
  wire [2:0] v_1478_0;
  wire [2:0] v_1479_0;
  wire [2:0] v_1480_0;
  reg [2:0] v_1481_0 = 3'h0;
  wire [0:0] v_1482_0;
  wire [0:0] v_1483_0;
  wire [0:0] v_1484_0;
  wire [2:0] v_1485_0;
  wire [2:0] v_1486_0;
  wire [2:0] v_1487_0;
  reg [2:0] v_1488_0 = 3'h0;
  wire [0:0] v_1489_0;
  wire [0:0] v_1490_0;
  wire [0:0] v_1491_0;
  wire [2:0] v_1492_0;
  wire [2:0] v_1493_0;
  wire [2:0] v_1494_0;
  reg [2:0] v_1495_0 = 3'h0;
  wire [0:0] v_1496_0;
  wire [0:0] v_1497_0;
  wire [0:0] v_1498_0;
  wire [2:0] v_1499_0;
  wire [2:0] v_1500_0;
  wire [2:0] v_1501_0;
  reg [2:0] v_1502_0 = 3'h0;
  wire [0:0] v_1503_0;
  wire [0:0] v_1504_0;
  wire [0:0] v_1505_0;
  wire [2:0] v_1506_0;
  wire [2:0] v_1507_0;
  wire [2:0] v_1508_0;
  reg [2:0] v_1509_0 = 3'h0;
  wire [0:0] v_1510_0;
  wire [0:0] v_1511_0;
  wire [0:0] v_1512_0;
  wire [2:0] v_1513_0;
  wire [2:0] v_1514_0;
  wire [2:0] v_1515_0;
  reg [2:0] v_1516_0 = 3'h0;
  wire [0:0] v_1517_0;
  wire [0:0] v_1518_0;
  wire [0:0] v_1519_0;
  wire [2:0] v_1520_0;
  wire [2:0] v_1521_0;
  wire [2:0] v_1522_0;
  reg [2:0] v_1523_0 = 3'h0;
  wire [0:0] v_1524_0;
  wire [0:0] v_1525_0;
  wire [0:0] v_1526_0;
  wire [2:0] v_1527_0;
  wire [2:0] v_1528_0;
  wire [2:0] v_1529_0;
  reg [2:0] v_1530_0 = 3'h0;
  wire [0:0] v_1531_0;
  wire [0:0] v_1532_0;
  wire [0:0] v_1533_0;
  wire [2:0] v_1534_0;
  wire [2:0] v_1535_0;
  wire [2:0] v_1536_0;
  reg [2:0] v_1537_0 = 3'h0;
  wire [0:0] v_1538_0;
  wire [0:0] v_1539_0;
  wire [0:0] v_1540_0;
  wire [2:0] v_1541_0;
  wire [2:0] v_1542_0;
  wire [2:0] v_1543_0;
  reg [2:0] v_1544_0 = 3'h0;
  wire [0:0] v_1545_0;
  wire [0:0] v_1546_0;
  wire [0:0] v_1547_0;
  wire [2:0] v_1548_0;
  wire [2:0] v_1549_0;
  wire [2:0] v_1550_0;
  reg [2:0] v_1551_0 = 3'h0;
  wire [0:0] v_1552_0;
  wire [0:0] v_1553_0;
  wire [0:0] v_1554_0;
  wire [2:0] v_1555_0;
  wire [2:0] v_1556_0;
  wire [2:0] v_1557_0;
  reg [2:0] v_1558_0 = 3'h0;
  wire [0:0] v_1559_0;
  wire [0:0] v_1560_0;
  wire [0:0] v_1561_0;
  wire [2:0] v_1562_0;
  wire [2:0] v_1563_0;
  wire [2:0] v_1564_0;
  reg [2:0] v_1565_0 = 3'h0;
  wire [0:0] v_1566_0;
  wire [0:0] v_1567_0;
  wire [0:0] v_1568_0;
  wire [2:0] v_1569_0;
  wire [2:0] v_1570_0;
  wire [2:0] v_1571_0;
  reg [2:0] v_1572_0 = 3'h0;
  wire [0:0] v_1573_0;
  wire [0:0] v_1574_0;
  wire [0:0] v_1575_0;
  wire [2:0] v_1576_0;
  wire [2:0] v_1577_0;
  wire [2:0] v_1578_0;
  reg [2:0] v_1579_0 = 3'h0;
  wire [0:0] v_1580_0;
  wire [0:0] v_1581_0;
  wire [0:0] v_1582_0;
  wire [2:0] v_1583_0;
  wire [2:0] v_1584_0;
  wire [2:0] v_1585_0;
  reg [2:0] v_1586_0 = 3'h0;
  wire [0:0] v_1587_0;
  wire [0:0] v_1588_0;
  wire [0:0] v_1589_0;
  wire [2:0] v_1590_0;
  wire [2:0] v_1591_0;
  wire [2:0] v_1592_0;
  reg [2:0] v_1593_0 = 3'h0;
  wire [0:0] v_1594_0;
  wire [0:0] v_1595_0;
  wire [0:0] v_1596_0;
  wire [2:0] v_1597_0;
  wire [2:0] v_1598_0;
  wire [2:0] v_1599_0;
  reg [2:0] v_1600_0 = 3'h0;
  wire [0:0] v_1601_0;
  wire [0:0] v_1602_0;
  wire [0:0] v_1603_0;
  wire [2:0] v_1604_0;
  wire [2:0] v_1605_0;
  wire [2:0] v_1606_0;
  reg [2:0] v_1607_0 = 3'h0;
  wire [0:0] v_1608_0;
  wire [0:0] v_1609_0;
  wire [0:0] v_1610_0;
  wire [2:0] v_1611_0;
  wire [2:0] v_1612_0;
  wire [2:0] v_1613_0;
  reg [2:0] v_1614_0 = 3'h0;
  wire [0:0] v_1615_0;
  wire [0:0] v_1616_0;
  wire [0:0] v_1617_0;
  wire [2:0] v_1618_0;
  wire [2:0] v_1619_0;
  wire [2:0] v_1620_0;
  reg [2:0] v_1621_0 = 3'h0;
  wire [0:0] v_1622_0;
  wire [0:0] v_1623_0;
  wire [0:0] v_1624_0;
  wire [2:0] v_1625_0;
  wire [2:0] v_1626_0;
  wire [2:0] v_1627_0;
  reg [2:0] v_1628_0 = 3'h0;
  wire [0:0] v_1629_0;
  wire [0:0] v_1630_0;
  wire [0:0] v_1631_0;
  wire [2:0] v_1632_0;
  wire [2:0] v_1633_0;
  wire [2:0] v_1634_0;
  reg [2:0] v_1635_0 = 3'h0;
  wire [0:0] v_1636_0;
  wire [0:0] v_1637_0;
  wire [0:0] v_1638_0;
  wire [2:0] v_1639_0;
  wire [2:0] v_1640_0;
  wire [2:0] v_1641_0;
  reg [2:0] v_1642_0 = 3'h0;
  wire [0:0] v_1643_0;
  wire [0:0] v_1644_0;
  wire [0:0] v_1645_0;
  wire [2:0] v_1646_0;
  wire [2:0] v_1647_0;
  wire [2:0] v_1648_0;
  reg [2:0] v_1649_0 = 3'h0;
  wire [0:0] v_1650_0;
  wire [0:0] v_1651_0;
  wire [0:0] v_1652_0;
  wire [2:0] v_1653_0;
  wire [2:0] v_1654_0;
  wire [2:0] v_1655_0;
  reg [2:0] v_1656_0 = 3'h0;
  wire [0:0] v_1657_0;
  wire [0:0] v_1658_0;
  wire [0:0] v_1659_0;
  wire [2:0] v_1660_0;
  wire [2:0] v_1661_0;
  wire [2:0] v_1662_0;
  reg [2:0] v_1663_0 = 3'h0;
  wire [0:0] v_1664_0;
  wire [0:0] v_1665_0;
  wire [0:0] v_1666_0;
  wire [2:0] v_1667_0;
  wire [2:0] v_1668_0;
  wire [2:0] v_1669_0;
  reg [2:0] v_1670_0 = 3'h0;
  wire [0:0] v_1671_0;
  wire [0:0] v_1672_0;
  wire [0:0] v_1673_0;
  wire [2:0] v_1674_0;
  wire [2:0] v_1675_0;
  wire [2:0] v_1676_0;
  reg [2:0] v_1677_0 = 3'h0;
  wire [0:0] v_1678_0;
  wire [0:0] v_1679_0;
  wire [0:0] v_1680_0;
  wire [2:0] v_1681_0;
  wire [2:0] v_1682_0;
  wire [2:0] v_1683_0;
  reg [2:0] v_1684_0 = 3'h0;
  wire [0:0] v_1685_0;
  wire [0:0] v_1686_0;
  wire [0:0] v_1687_0;
  wire [2:0] v_1688_0;
  wire [2:0] v_1689_0;
  wire [2:0] v_1690_0;
  reg [2:0] v_1691_0 = 3'h0;
  wire [0:0] v_1692_0;
  wire [0:0] v_1693_0;
  wire [0:0] v_1694_0;
  wire [2:0] v_1695_0;
  wire [2:0] v_1696_0;
  wire [2:0] v_1697_0;
  reg [2:0] v_1698_0 = 3'h0;
  wire [0:0] v_1699_0;
  wire [0:0] v_1700_0;
  wire [0:0] v_1701_0;
  wire [2:0] v_1702_0;
  wire [2:0] v_1703_0;
  wire [2:0] v_1704_0;
  reg [2:0] v_1705_0 = 3'h0;
  wire [0:0] v_1706_0;
  wire [0:0] v_1707_0;
  wire [0:0] v_1708_0;
  wire [2:0] v_1709_0;
  wire [2:0] v_1710_0;
  wire [2:0] v_1711_0;
  reg [2:0] v_1712_0 = 3'h0;
  wire [0:0] v_1713_0;
  wire [0:0] v_1714_0;
  wire [0:0] v_1715_0;
  wire [2:0] v_1716_0;
  wire [2:0] v_1717_0;
  wire [2:0] v_1718_0;
  reg [2:0] v_1719_0 = 3'h0;
  wire [0:0] v_1720_0;
  wire [0:0] v_1721_0;
  wire [0:0] v_1722_0;
  wire [2:0] v_1723_0;
  wire [2:0] v_1724_0;
  wire [2:0] v_1725_0;
  reg [2:0] v_1726_0 = 3'h0;
  wire [0:0] v_1727_0;
  wire [0:0] v_1728_0;
  wire [0:0] v_1729_0;
  wire [2:0] v_1730_0;
  wire [2:0] v_1731_0;
  wire [2:0] v_1732_0;
  reg [2:0] v_1733_0 = 3'h0;
  wire [0:0] v_1734_0;
  wire [0:0] v_1735_0;
  wire [0:0] v_1736_0;
  wire [2:0] v_1737_0;
  wire [2:0] v_1738_0;
  wire [2:0] v_1739_0;
  reg [2:0] v_1740_0 = 3'h0;
  wire [0:0] v_1741_0;
  wire [0:0] v_1742_0;
  wire [0:0] v_1743_0;
  wire [2:0] v_1744_0;
  wire [2:0] v_1745_0;
  wire [2:0] v_1746_0;
  reg [2:0] v_1747_0 = 3'h0;
  wire [0:0] v_1748_0;
  wire [0:0] v_1749_0;
  wire [0:0] v_1750_0;
  wire [2:0] v_1751_0;
  wire [2:0] v_1752_0;
  wire [2:0] v_1753_0;
  reg [2:0] v_1754_0 = 3'h0;
  wire [0:0] v_1755_0;
  wire [0:0] v_1756_0;
  wire [0:0] v_1757_0;
  wire [2:0] v_1758_0;
  wire [2:0] v_1759_0;
  wire [2:0] v_1760_0;
  reg [2:0] v_1761_0 = 3'h0;
  wire [0:0] v_1762_0;
  wire [0:0] v_1763_0;
  wire [0:0] v_1764_0;
  wire [2:0] v_1765_0;
  wire [2:0] v_1766_0;
  wire [2:0] v_1767_0;
  reg [2:0] v_1768_0 = 3'h0;
  wire [0:0] v_1769_0;
  wire [0:0] v_1770_0;
  wire [0:0] v_1771_0;
  wire [2:0] v_1772_0;
  wire [2:0] v_1773_0;
  wire [2:0] v_1774_0;
  reg [2:0] v_1775_0 = 3'h0;
  wire [0:0] v_1776_0;
  wire [0:0] v_1777_0;
  wire [0:0] v_1778_0;
  wire [2:0] v_1779_0;
  wire [2:0] v_1780_0;
  wire [2:0] v_1781_0;
  reg [2:0] v_1782_0 = 3'h0;
  wire [0:0] v_1783_0;
  wire [0:0] v_1784_0;
  wire [0:0] v_1785_0;
  wire [2:0] v_1786_0;
  wire [2:0] v_1787_0;
  wire [2:0] v_1788_0;
  reg [2:0] v_1789_0 = 3'h0;
  wire [0:0] v_1790_0;
  wire [0:0] v_1791_0;
  wire [0:0] v_1792_0;
  wire [2:0] v_1793_0;
  wire [2:0] v_1794_0;
  wire [2:0] v_1795_0;
  reg [2:0] v_1796_0 = 3'h0;
  wire [0:0] v_1797_0;
  wire [0:0] v_1798_0;
  wire [0:0] v_1799_0;
  wire [2:0] v_1800_0;
  wire [2:0] v_1801_0;
  wire [2:0] v_1802_0;
  reg [2:0] v_1803_0 = 3'h0;
  wire [0:0] v_1804_0;
  wire [0:0] v_1805_0;
  wire [0:0] v_1806_0;
  wire [2:0] v_1807_0;
  wire [2:0] v_1808_0;
  wire [2:0] v_1809_0;
  reg [2:0] v_1810_0 = 3'h0;
  wire [0:0] v_1811_0;
  wire [0:0] v_1812_0;
  wire [0:0] v_1813_0;
  wire [2:0] v_1814_0;
  wire [2:0] v_1815_0;
  wire [2:0] v_1816_0;
  reg [2:0] v_1817_0 = 3'h0;
  wire [0:0] v_1818_0;
  wire [0:0] v_1819_0;
  wire [0:0] v_1820_0;
  wire [2:0] v_1821_0;
  wire [2:0] v_1822_0;
  wire [2:0] v_1823_0;
  reg [2:0] v_1824_0 = 3'h0;
  wire [0:0] v_1825_0;
  wire [0:0] v_1826_0;
  wire [0:0] v_1827_0;
  wire [2:0] v_1828_0;
  wire [2:0] v_1829_0;
  wire [2:0] v_1830_0;
  reg [2:0] v_1831_0 = 3'h0;
  wire [0:0] v_1832_0;
  wire [0:0] v_1833_0;
  wire [0:0] v_1834_0;
  wire [2:0] v_1835_0;
  wire [2:0] v_1836_0;
  wire [2:0] v_1837_0;
  reg [2:0] v_1838_0 = 3'h0;
  wire [0:0] v_1839_0;
  wire [0:0] v_1840_0;
  wire [0:0] v_1841_0;
  wire [2:0] v_1842_0;
  wire [2:0] v_1843_0;
  wire [2:0] v_1844_0;
  reg [2:0] v_1845_0 = 3'h0;
  wire [0:0] v_1846_0;
  wire [0:0] v_1847_0;
  wire [0:0] v_1848_0;
  wire [2:0] v_1849_0;
  wire [2:0] v_1850_0;
  wire [2:0] v_1851_0;
  reg [2:0] v_1852_0 = 3'h0;
  wire [0:0] v_1853_0;
  wire [0:0] v_1854_0;
  wire [0:0] v_1855_0;
  wire [2:0] v_1856_0;
  wire [2:0] v_1857_0;
  wire [2:0] v_1858_0;
  reg [2:0] v_1859_0 = 3'h0;
  wire [0:0] v_1860_0;
  wire [0:0] v_1861_0;
  wire [0:0] v_1862_0;
  wire [2:0] v_1863_0;
  wire [2:0] v_1864_0;
  wire [2:0] v_1865_0;
  reg [2:0] v_1866_0 = 3'h0;
  wire [0:0] v_1867_0;
  wire [0:0] v_1868_0;
  wire [0:0] v_1869_0;
  wire [2:0] v_1870_0;
  wire [2:0] v_1871_0;
  wire [2:0] v_1872_0;
  reg [2:0] v_1873_0 = 3'h0;
  wire [0:0] v_1874_0;
  wire [0:0] v_1875_0;
  wire [0:0] v_1876_0;
  wire [2:0] v_1877_0;
  wire [2:0] v_1878_0;
  wire [2:0] v_1879_0;
  reg [2:0] v_1880_0 = 3'h0;
  wire [0:0] v_1881_0;
  wire [0:0] v_1882_0;
  wire [0:0] v_1883_0;
  wire [2:0] v_1884_0;
  wire [2:0] v_1885_0;
  wire [2:0] v_1886_0;
  reg [2:0] v_1887_0 = 3'h0;
  wire [0:0] v_1888_0;
  wire [0:0] v_1889_0;
  wire [0:0] v_1890_0;
  wire [2:0] v_1891_0;
  wire [2:0] v_1892_0;
  wire [2:0] v_1893_0;
  reg [2:0] v_1894_0 = 3'h0;
  wire [0:0] v_1895_0;
  wire [0:0] v_1896_0;
  wire [0:0] v_1897_0;
  wire [2:0] v_1898_0;
  wire [2:0] v_1899_0;
  wire [2:0] v_1900_0;
  reg [2:0] v_1901_0 = 3'h0;
  wire [0:0] v_1902_0;
  wire [0:0] v_1903_0;
  wire [0:0] v_1904_0;
  wire [2:0] v_1905_0;
  wire [2:0] v_1906_0;
  wire [2:0] v_1907_0;
  reg [2:0] v_1908_0 = 3'h0;
  wire [0:0] v_1909_0;
  wire [0:0] v_1910_0;
  wire [0:0] v_1911_0;
  wire [2:0] v_1912_0;
  wire [2:0] v_1913_0;
  wire [2:0] v_1914_0;
  reg [2:0] v_1915_0 = 3'h0;
  wire [0:0] v_1916_0;
  wire [0:0] v_1917_0;
  wire [0:0] v_1918_0;
  wire [2:0] v_1919_0;
  wire [2:0] v_1920_0;
  wire [2:0] v_1921_0;
  reg [2:0] v_1922_0 = 3'h0;
  wire [0:0] v_1923_0;
  wire [0:0] v_1924_0;
  wire [0:0] v_1925_0;
  wire [2:0] v_1926_0;
  wire [2:0] v_1927_0;
  wire [2:0] v_1928_0;
  reg [2:0] v_1929_0 = 3'h0;
  wire [0:0] v_1930_0;
  wire [0:0] v_1931_0;
  wire [0:0] v_1932_0;
  wire [2:0] v_1933_0;
  wire [2:0] v_1934_0;
  wire [2:0] v_1935_0;
  reg [2:0] v_1936_0 = 3'h0;
  wire [0:0] v_1937_0;
  wire [0:0] v_1938_0;
  wire [0:0] v_1939_0;
  wire [2:0] v_1940_0;
  wire [2:0] v_1941_0;
  wire [2:0] v_1942_0;
  reg [2:0] v_1943_0 = 3'h0;
  wire [0:0] v_1944_0;
  wire [0:0] v_1945_0;
  wire [0:0] v_1946_0;
  wire [2:0] v_1947_0;
  wire [2:0] v_1948_0;
  wire [2:0] v_1949_0;
  reg [2:0] v_1950_0 = 3'h0;
  wire [0:0] v_1951_0;
  wire [0:0] v_1952_0;
  wire [0:0] v_1953_0;
  wire [2:0] v_1954_0;
  wire [2:0] v_1955_0;
  wire [2:0] v_1956_0;
  reg [2:0] v_1957_0 = 3'h0;
  wire [0:0] v_1958_0;
  wire [0:0] v_1959_0;
  wire [0:0] v_1960_0;
  wire [2:0] v_1961_0;
  wire [2:0] v_1962_0;
  wire [2:0] v_1963_0;
  reg [2:0] v_1964_0 = 3'h0;
  wire [0:0] v_1965_0;
  wire [0:0] v_1966_0;
  wire [0:0] v_1967_0;
  wire [2:0] v_1968_0;
  wire [2:0] v_1969_0;
  wire [2:0] v_1970_0;
  reg [2:0] v_1971_0 = 3'h0;
  wire [0:0] v_1972_0;
  wire [0:0] v_1973_0;
  wire [0:0] v_1974_0;
  wire [2:0] v_1975_0;
  wire [2:0] v_1976_0;
  wire [2:0] v_1977_0;
  reg [2:0] v_1978_0 = 3'h0;
  wire [0:0] v_1979_0;
  wire [0:0] v_1980_0;
  wire [0:0] v_1981_0;
  wire [2:0] v_1982_0;
  wire [2:0] v_1983_0;
  wire [2:0] v_1984_0;
  reg [2:0] v_1985_0 = 3'h0;
  wire [0:0] v_1986_0;
  wire [0:0] v_1987_0;
  wire [0:0] v_1988_0;
  wire [2:0] v_1989_0;
  wire [2:0] v_1990_0;
  wire [2:0] v_1991_0;
  reg [2:0] v_1992_0 = 3'h0;
  wire [0:0] v_1993_0;
  wire [0:0] v_1994_0;
  wire [0:0] v_1995_0;
  wire [2:0] v_1996_0;
  wire [2:0] v_1997_0;
  wire [2:0] v_1998_0;
  reg [2:0] v_1999_0 = 3'h0;
  wire [0:0] v_2000_0;
  wire [0:0] v_2001_0;
  wire [0:0] v_2002_0;
  wire [2:0] v_2003_0;
  wire [2:0] v_2004_0;
  wire [2:0] v_2005_0;
  reg [2:0] v_2006_0 = 3'h0;
  wire [0:0] v_2007_0;
  wire [0:0] v_2008_0;
  wire [0:0] v_2009_0;
  wire [2:0] v_2010_0;
  wire [2:0] v_2011_0;
  wire [2:0] v_2012_0;
  reg [2:0] v_2013_0 = 3'h0;
  wire [0:0] v_2014_0;
  wire [0:0] v_2015_0;
  wire [0:0] v_2016_0;
  wire [2:0] v_2017_0;
  wire [2:0] v_2018_0;
  wire [2:0] v_2019_0;
  reg [2:0] v_2020_0 = 3'h0;
  wire [0:0] v_2021_0;
  wire [0:0] v_2022_0;
  wire [0:0] v_2023_0;
  wire [2:0] v_2024_0;
  wire [2:0] v_2025_0;
  wire [2:0] v_2026_0;
  reg [2:0] v_2027_0 = 3'h0;
  wire [0:0] v_2028_0;
  wire [0:0] v_2029_0;
  wire [0:0] v_2030_0;
  wire [2:0] v_2031_0;
  wire [2:0] v_2032_0;
  wire [2:0] v_2033_0;
  reg [2:0] v_2034_0 = 3'h0;
  wire [0:0] v_2035_0;
  wire [0:0] v_2036_0;
  wire [0:0] v_2037_0;
  wire [2:0] v_2038_0;
  wire [2:0] v_2039_0;
  wire [2:0] v_2040_0;
  reg [2:0] v_2041_0 = 3'h0;
  wire [0:0] v_2042_0;
  wire [0:0] v_2043_0;
  wire [0:0] v_2044_0;
  wire [2:0] v_2045_0;
  wire [2:0] v_2046_0;
  wire [2:0] v_2047_0;
  reg [2:0] v_2048_0 = 3'h0;
  wire [0:0] v_2049_0;
  wire [0:0] v_2050_0;
  wire [0:0] v_2051_0;
  wire [2:0] v_2052_0;
  wire [2:0] v_2053_0;
  wire [2:0] v_2054_0;
  reg [2:0] v_2055_0 = 3'h0;
  wire [0:0] v_2056_0;
  wire [0:0] v_2057_0;
  wire [0:0] v_2058_0;
  wire [2:0] v_2059_0;
  wire [2:0] v_2060_0;
  wire [2:0] v_2061_0;
  reg [2:0] v_2062_0 = 3'h0;
  wire [0:0] v_2063_0;
  wire [0:0] v_2064_0;
  wire [0:0] v_2065_0;
  wire [2:0] v_2066_0;
  wire [2:0] v_2067_0;
  wire [2:0] v_2068_0;
  reg [2:0] v_2069_0 = 3'h0;
  wire [0:0] v_2070_0;
  wire [0:0] v_2071_0;
  wire [0:0] v_2072_0;
  wire [2:0] v_2073_0;
  wire [2:0] v_2074_0;
  wire [2:0] v_2075_0;
  reg [2:0] v_2076_0 = 3'h0;
  wire [0:0] v_2077_0;
  wire [0:0] v_2078_0;
  wire [0:0] v_2079_0;
  wire [2:0] v_2080_0;
  wire [2:0] v_2081_0;
  wire [2:0] v_2082_0;
  reg [2:0] v_2083_0 = 3'h0;
  wire [0:0] v_2084_0;
  wire [0:0] v_2085_0;
  wire [0:0] v_2086_0;
  wire [2:0] v_2087_0;
  wire [2:0] v_2088_0;
  wire [2:0] v_2089_0;
  reg [2:0] v_2090_0 = 3'h0;
  wire [0:0] v_2091_0;
  wire [0:0] v_2092_0;
  wire [0:0] v_2093_0;
  wire [2:0] v_2094_0;
  wire [2:0] v_2095_0;
  wire [2:0] v_2096_0;
  reg [2:0] v_2097_0 = 3'h0;
  wire [0:0] v_2098_0;
  wire [0:0] v_2099_0;
  wire [0:0] v_2100_0;
  wire [2:0] v_2101_0;
  wire [2:0] v_2102_0;
  wire [2:0] v_2103_0;
  reg [2:0] v_2104_0 = 3'h0;
  wire [0:0] v_2105_0;
  wire [0:0] v_2106_0;
  wire [0:0] v_2107_0;
  wire [2:0] v_2108_0;
  wire [2:0] v_2109_0;
  wire [2:0] v_2110_0;
  reg [2:0] v_2111_0 = 3'h0;
  wire [0:0] v_2112_0;
  wire [0:0] v_2113_0;
  wire [0:0] v_2114_0;
  wire [2:0] v_2115_0;
  wire [2:0] v_2116_0;
  wire [2:0] v_2117_0;
  reg [2:0] v_2118_0 = 3'h0;
  wire [0:0] v_2119_0;
  wire [0:0] v_2120_0;
  wire [0:0] v_2121_0;
  wire [2:0] v_2122_0;
  wire [2:0] v_2123_0;
  wire [2:0] v_2124_0;
  reg [2:0] v_2125_0 = 3'h0;
  wire [0:0] v_2126_0;
  wire [0:0] v_2127_0;
  wire [0:0] v_2128_0;
  wire [2:0] v_2129_0;
  wire [2:0] v_2130_0;
  wire [2:0] v_2131_0;
  reg [2:0] v_2132_0 = 3'h0;
  wire [0:0] v_2133_0;
  wire [0:0] v_2134_0;
  wire [0:0] v_2135_0;
  wire [2:0] v_2136_0;
  wire [2:0] v_2137_0;
  wire [2:0] v_2138_0;
  reg [2:0] v_2139_0 = 3'h0;
  wire [0:0] v_2140_0;
  wire [0:0] v_2141_0;
  wire [0:0] v_2142_0;
  wire [2:0] v_2143_0;
  wire [2:0] v_2144_0;
  wire [2:0] v_2145_0;
  reg [2:0] v_2146_0 = 3'h0;
  wire [0:0] v_2147_0;
  wire [0:0] v_2148_0;
  wire [0:0] v_2149_0;
  wire [2:0] v_2150_0;
  wire [2:0] v_2151_0;
  wire [2:0] v_2152_0;
  reg [2:0] v_2153_0 = 3'h0;
  wire [0:0] v_2154_0;
  wire [0:0] v_2155_0;
  wire [0:0] v_2156_0;
  wire [2:0] v_2157_0;
  wire [2:0] v_2158_0;
  wire [2:0] v_2159_0;
  reg [2:0] v_2160_0 = 3'h0;
  wire [0:0] v_2161_0;
  wire [0:0] v_2162_0;
  wire [0:0] v_2163_0;
  wire [2:0] v_2164_0;
  wire [2:0] v_2165_0;
  wire [2:0] v_2166_0;
  reg [2:0] v_2167_0 = 3'h0;
  wire [0:0] v_2168_0;
  wire [0:0] v_2169_0;
  wire [0:0] v_2170_0;
  wire [2:0] v_2171_0;
  wire [2:0] v_2172_0;
  wire [2:0] v_2173_0;
  reg [2:0] v_2174_0 = 3'h0;
  wire [0:0] v_2175_0;
  wire [0:0] v_2176_0;
  wire [0:0] v_2177_0;
  wire [2:0] v_2178_0;
  wire [2:0] v_2179_0;
  wire [2:0] v_2180_0;
  reg [2:0] v_2181_0 = 3'h0;
  wire [0:0] v_2182_0;
  wire [0:0] v_2183_0;
  wire [0:0] v_2184_0;
  wire [2:0] v_2185_0;
  wire [2:0] v_2186_0;
  wire [2:0] v_2187_0;
  reg [2:0] v_2188_0 = 3'h0;
  wire [0:0] v_2189_0;
  wire [0:0] v_2190_0;
  wire [0:0] v_2191_0;
  wire [2:0] v_2192_0;
  wire [2:0] v_2193_0;
  wire [2:0] v_2194_0;
  reg [2:0] v_2195_0 = 3'h0;
  wire [0:0] v_2196_0;
  wire [0:0] v_2197_0;
  wire [0:0] v_2198_0;
  wire [2:0] v_2199_0;
  wire [2:0] v_2200_0;
  wire [2:0] v_2201_0;
  reg [2:0] v_2202_0 = 3'h0;
  wire [0:0] v_2203_0;
  wire [0:0] v_2204_0;
  wire [0:0] v_2205_0;
  wire [2:0] v_2206_0;
  wire [2:0] v_2207_0;
  wire [2:0] v_2208_0;
  reg [2:0] v_2209_0 = 3'h0;
  wire [0:0] v_2210_0;
  wire [0:0] v_2211_0;
  wire [0:0] v_2212_0;
  wire [2:0] v_2213_0;
  wire [2:0] v_2214_0;
  wire [2:0] v_2215_0;
  reg [2:0] v_2216_0 = 3'h0;
  wire [0:0] v_2217_0;
  wire [0:0] v_2218_0;
  wire [0:0] v_2219_0;
  wire [2:0] v_2220_0;
  wire [2:0] v_2221_0;
  wire [2:0] v_2222_0;
  reg [2:0] v_2223_0 = 3'h0;
  wire [0:0] v_2224_0;
  wire [0:0] v_2225_0;
  wire [0:0] v_2226_0;
  wire [2:0] v_2227_0;
  wire [2:0] v_2228_0;
  wire [2:0] v_2229_0;
  reg [2:0] v_2230_0 = 3'h0;
  wire [0:0] v_2231_0;
  wire [0:0] v_2232_0;
  wire [0:0] v_2233_0;
  wire [2:0] v_2234_0;
  wire [2:0] v_2235_0;
  wire [2:0] v_2236_0;
  reg [2:0] v_2237_0 = 3'h0;
  wire [0:0] v_2238_0;
  wire [0:0] v_2239_0;
  wire [0:0] v_2240_0;
  wire [2:0] v_2241_0;
  wire [2:0] v_2242_0;
  wire [2:0] v_2243_0;
  reg [2:0] v_2244_0 = 3'h0;
  wire [0:0] v_2245_0;
  wire [0:0] v_2246_0;
  wire [0:0] v_2247_0;
  wire [2:0] v_2248_0;
  wire [2:0] v_2249_0;
  wire [2:0] v_2250_0;
  reg [2:0] v_2251_0 = 3'h0;
  wire [0:0] v_2252_0;
  wire [0:0] v_2253_0;
  wire [0:0] v_2254_0;
  wire [2:0] v_2255_0;
  wire [2:0] v_2256_0;
  wire [2:0] v_2257_0;
  reg [2:0] v_2258_0 = 3'h0;
  wire [0:0] v_2259_0;
  wire [0:0] v_2260_0;
  wire [0:0] v_2261_0;
  wire [2:0] v_2262_0;
  wire [2:0] v_2263_0;
  wire [2:0] v_2264_0;
  reg [2:0] v_2265_0 = 3'h0;
  wire [0:0] v_2266_0;
  wire [0:0] v_2267_0;
  wire [0:0] v_2268_0;
  wire [2:0] v_2269_0;
  wire [2:0] v_2270_0;
  wire [2:0] v_2271_0;
  reg [2:0] v_2272_0 = 3'h0;
  wire [0:0] v_2273_0;
  wire [0:0] v_2274_0;
  wire [0:0] v_2275_0;
  wire [2:0] v_2276_0;
  wire [2:0] v_2277_0;
  wire [2:0] v_2278_0;
  reg [2:0] v_2279_0 = 3'h0;
  wire [0:0] v_2280_0;
  wire [0:0] v_2281_0;
  wire [0:0] v_2282_0;
  wire [2:0] v_2283_0;
  wire [2:0] v_2284_0;
  wire [2:0] v_2285_0;
  reg [2:0] v_2286_0 = 3'h0;
  wire [0:0] v_2287_0;
  wire [0:0] v_2288_0;
  wire [0:0] v_2289_0;
  wire [2:0] v_2290_0;
  wire [2:0] v_2291_0;
  wire [2:0] v_2292_0;
  reg [2:0] v_2293_0 = 3'h0;
  wire [0:0] v_2294_0;
  wire [0:0] v_2295_0;
  wire [0:0] v_2296_0;
  wire [2:0] v_2297_0;
  wire [2:0] v_2298_0;
  wire [2:0] v_2299_0;
  reg [2:0] v_2300_0 = 3'h0;
  wire [0:0] v_2301_0;
  wire [0:0] v_2302_0;
  wire [0:0] v_2303_0;
  wire [2:0] v_2304_0;
  wire [2:0] v_2305_0;
  wire [2:0] v_2306_0;
  reg [2:0] v_2307_0 = 3'h0;
  wire [0:0] v_2308_0;
  wire [0:0] v_2309_0;
  wire [0:0] v_2310_0;
  wire [2:0] v_2311_0;
  wire [2:0] v_2312_0;
  wire [2:0] v_2313_0;
  reg [2:0] v_2314_0 = 3'h0;
  wire [0:0] v_2315_0;
  wire [0:0] v_2316_0;
  wire [0:0] v_2317_0;
  wire [2:0] v_2318_0;
  wire [2:0] v_2319_0;
  wire [2:0] v_2320_0;
  reg [2:0] v_2321_0 = 3'h0;
  wire [0:0] v_2322_0;
  wire [0:0] v_2323_0;
  wire [0:0] v_2324_0;
  wire [2:0] v_2325_0;
  wire [2:0] v_2326_0;
  wire [2:0] v_2327_0;
  reg [2:0] v_2328_0 = 3'h0;
  wire [0:0] v_2329_0;
  wire [0:0] v_2330_0;
  wire [0:0] v_2331_0;
  wire [2:0] v_2332_0;
  wire [2:0] v_2333_0;
  wire [2:0] v_2334_0;
  reg [2:0] v_2335_0 = 3'h0;
  wire [0:0] v_2336_0;
  wire [0:0] v_2337_0;
  wire [0:0] v_2338_0;
  wire [2:0] v_2339_0;
  wire [2:0] v_2340_0;
  wire [2:0] v_2341_0;
  reg [2:0] v_2342_0 = 3'h0;
  wire [0:0] v_2343_0;
  wire [0:0] v_2344_0;
  wire [0:0] v_2345_0;
  wire [2:0] v_2346_0;
  wire [2:0] v_2347_0;
  wire [2:0] v_2348_0;
  reg [2:0] v_2349_0 = 3'h0;
  wire [0:0] v_2350_0;
  wire [0:0] v_2351_0;
  wire [0:0] v_2352_0;
  wire [2:0] v_2353_0;
  wire [2:0] v_2354_0;
  wire [2:0] v_2355_0;
  reg [2:0] v_2356_0 = 3'h0;
  wire [0:0] v_2357_0;
  wire [0:0] v_2358_0;
  wire [0:0] v_2359_0;
  wire [2:0] v_2360_0;
  wire [2:0] v_2361_0;
  wire [2:0] v_2362_0;
  reg [2:0] v_2363_0 = 3'h0;
  wire [0:0] v_2364_0;
  wire [0:0] v_2365_0;
  wire [0:0] v_2366_0;
  wire [2:0] v_2367_0;
  wire [2:0] v_2368_0;
  wire [2:0] v_2369_0;
  reg [2:0] v_2370_0 = 3'h0;
  wire [0:0] v_2371_0;
  wire [0:0] v_2372_0;
  wire [0:0] v_2373_0;
  wire [2:0] v_2374_0;
  wire [2:0] v_2375_0;
  wire [2:0] v_2376_0;
  reg [2:0] v_2377_0 = 3'h0;
  wire [0:0] v_2378_0;
  wire [0:0] v_2379_0;
  wire [0:0] v_2380_0;
  wire [2:0] v_2381_0;
  wire [2:0] v_2382_0;
  wire [2:0] v_2383_0;
  reg [2:0] v_2384_0 = 3'h0;
  wire [0:0] v_2385_0;
  wire [0:0] v_2386_0;
  wire [0:0] v_2387_0;
  wire [2:0] v_2388_0;
  wire [2:0] v_2389_0;
  wire [2:0] v_2390_0;
  reg [2:0] v_2391_0 = 3'h0;
  wire [0:0] v_2392_0;
  wire [0:0] v_2393_0;
  wire [0:0] v_2394_0;
  wire [2:0] v_2395_0;
  wire [2:0] v_2396_0;
  wire [2:0] v_2397_0;
  reg [2:0] v_2398_0 = 3'h0;
  wire [0:0] v_2399_0;
  wire [0:0] v_2400_0;
  wire [0:0] v_2401_0;
  wire [2:0] v_2402_0;
  wire [2:0] v_2403_0;
  wire [2:0] v_2404_0;
  reg [2:0] v_2405_0 = 3'h0;
  wire [0:0] v_2406_0;
  wire [0:0] v_2407_0;
  wire [0:0] v_2408_0;
  wire [2:0] v_2409_0;
  wire [2:0] v_2410_0;
  wire [2:0] v_2411_0;
  reg [2:0] v_2412_0 = 3'h0;
  wire [0:0] v_2413_0;
  wire [0:0] v_2414_0;
  wire [0:0] v_2415_0;
  wire [2:0] v_2416_0;
  wire [2:0] v_2417_0;
  wire [2:0] v_2418_0;
  reg [2:0] v_2419_0 = 3'h0;
  wire [0:0] v_2420_0;
  wire [0:0] v_2421_0;
  wire [0:0] v_2422_0;
  wire [2:0] v_2423_0;
  wire [2:0] v_2424_0;
  wire [2:0] v_2425_0;
  reg [2:0] v_2426_0 = 3'h0;
  wire [0:0] v_2427_0;
  wire [0:0] v_2428_0;
  wire [0:0] v_2429_0;
  wire [2:0] v_2430_0;
  wire [2:0] v_2431_0;
  wire [2:0] v_2432_0;
  reg [2:0] v_2433_0 = 3'h0;
  wire [0:0] v_2434_0;
  wire [0:0] v_2435_0;
  wire [0:0] v_2436_0;
  wire [2:0] v_2437_0;
  wire [2:0] v_2438_0;
  wire [2:0] v_2439_0;
  reg [2:0] v_2440_0 = 3'h0;
  wire [0:0] v_2441_0;
  wire [0:0] v_2442_0;
  wire [0:0] v_2443_0;
  wire [2:0] v_2444_0;
  wire [2:0] v_2445_0;
  wire [2:0] v_2446_0;
  reg [2:0] v_2447_0 = 3'h0;
  wire [0:0] v_2448_0;
  wire [0:0] v_2449_0;
  wire [0:0] v_2450_0;
  wire [2:0] v_2451_0;
  wire [2:0] v_2452_0;
  wire [2:0] v_2453_0;
  reg [2:0] v_2454_0 = 3'h0;
  wire [0:0] v_2455_0;
  wire [0:0] v_2456_0;
  wire [0:0] v_2457_0;
  wire [2:0] v_2458_0;
  wire [2:0] v_2459_0;
  wire [2:0] v_2460_0;
  reg [2:0] v_2461_0 = 3'h0;
  wire [0:0] v_2462_0;
  wire [0:0] v_2463_0;
  wire [0:0] v_2464_0;
  wire [2:0] v_2465_0;
  wire [2:0] v_2466_0;
  wire [2:0] v_2467_0;
  reg [2:0] v_2468_0 = 3'h0;
  wire [0:0] v_2469_0;
  wire [0:0] v_2470_0;
  wire [0:0] v_2471_0;
  wire [2:0] v_2472_0;
  wire [2:0] v_2473_0;
  wire [2:0] v_2474_0;
  reg [2:0] v_2475_0 = 3'h0;
  wire [0:0] v_2476_0;
  wire [0:0] v_2477_0;
  wire [0:0] v_2478_0;
  wire [2:0] v_2479_0;
  wire [2:0] v_2480_0;
  wire [2:0] v_2481_0;
  reg [2:0] v_2482_0 = 3'h0;
  wire [0:0] v_2483_0;
  wire [0:0] v_2484_0;
  wire [0:0] v_2485_0;
  wire [2:0] v_2486_0;
  wire [2:0] v_2487_0;
  wire [2:0] v_2488_0;
  reg [2:0] v_2489_0 = 3'h0;
  wire [0:0] v_2490_0;
  wire [0:0] v_2491_0;
  wire [0:0] v_2492_0;
  wire [2:0] v_2493_0;
  wire [2:0] v_2494_0;
  wire [2:0] v_2495_0;
  reg [2:0] v_2496_0 = 3'h0;
  wire [0:0] v_2497_0;
  wire [0:0] v_2498_0;
  wire [0:0] v_2499_0;
  wire [2:0] v_2500_0;
  wire [2:0] v_2501_0;
  wire [2:0] v_2502_0;
  reg [2:0] v_2503_0 = 3'h0;
  wire [0:0] v_2504_0;
  wire [0:0] v_2505_0;
  wire [0:0] v_2506_0;
  wire [2:0] v_2507_0;
  wire [2:0] v_2508_0;
  wire [2:0] v_2509_0;
  reg [2:0] v_2510_0 = 3'h0;
  wire [0:0] v_2511_0;
  wire [0:0] v_2512_0;
  wire [0:0] v_2513_0;
  wire [2:0] v_2514_0;
  wire [2:0] v_2515_0;
  wire [2:0] v_2516_0;
  reg [2:0] v_2517_0 = 3'h0;
  wire [0:0] v_2518_0;
  wire [0:0] v_2519_0;
  wire [0:0] v_2520_0;
  wire [2:0] v_2521_0;
  wire [2:0] v_2522_0;
  wire [2:0] v_2523_0;
  reg [2:0] v_2524_0 = 3'h0;
  wire [0:0] v_2525_0;
  wire [0:0] v_2526_0;
  wire [0:0] v_2527_0;
  wire [2:0] v_2528_0;
  wire [2:0] v_2529_0;
  wire [2:0] v_2530_0;
  reg [2:0] v_2531_0 = 3'h0;
  wire [0:0] v_2532_0;
  wire [0:0] v_2533_0;
  wire [0:0] v_2534_0;
  wire [2:0] v_2535_0;
  wire [2:0] v_2536_0;
  wire [2:0] v_2537_0;
  reg [2:0] v_2538_0 = 3'h0;
  wire [0:0] v_2539_0;
  wire [0:0] v_2540_0;
  wire [0:0] v_2541_0;
  wire [2:0] v_2542_0;
  wire [2:0] v_2543_0;
  wire [2:0] v_2544_0;
  reg [2:0] v_2545_0 = 3'h0;
  wire [0:0] v_2546_0;
  wire [0:0] v_2547_0;
  wire [0:0] v_2548_0;
  wire [2:0] v_2549_0;
  wire [2:0] v_2550_0;
  wire [2:0] v_2551_0;
  reg [2:0] v_2552_0 = 3'h0;
  wire [0:0] v_2553_0;
  wire [0:0] v_2554_0;
  wire [0:0] v_2555_0;
  wire [2:0] v_2556_0;
  wire [2:0] v_2557_0;
  wire [2:0] v_2558_0;
  reg [2:0] v_2559_0 = 3'h0;
  wire [0:0] v_2560_0;
  wire [0:0] v_2561_0;
  wire [0:0] v_2562_0;
  wire [2:0] v_2563_0;
  wire [2:0] v_2564_0;
  wire [2:0] v_2565_0;
  reg [2:0] v_2566_0 = 3'h0;
  wire [0:0] v_2567_0;
  wire [0:0] v_2568_0;
  wire [0:0] v_2569_0;
  wire [2:0] v_2570_0;
  wire [2:0] v_2571_0;
  wire [2:0] v_2572_0;
  reg [2:0] v_2573_0 = 3'h0;
  wire [0:0] v_2574_0;
  wire [0:0] v_2575_0;
  wire [0:0] v_2576_0;
  wire [2:0] v_2577_0;
  wire [2:0] v_2578_0;
  wire [2:0] v_2579_0;
  reg [2:0] v_2580_0 = 3'h0;
  wire [0:0] v_2581_0;
  wire [0:0] v_2582_0;
  wire [0:0] v_2583_0;
  wire [2:0] v_2584_0;
  wire [2:0] v_2585_0;
  wire [2:0] v_2586_0;
  reg [2:0] v_2587_0 = 3'h0;
  wire [0:0] v_2588_0;
  wire [0:0] v_2589_0;
  wire [0:0] v_2590_0;
  wire [2:0] v_2591_0;
  wire [2:0] v_2592_0;
  wire [2:0] v_2593_0;
  reg [2:0] v_2594_0 = 3'h0;
  wire [0:0] v_2595_0;
  wire [0:0] v_2596_0;
  wire [0:0] v_2597_0;
  wire [2:0] v_2598_0;
  wire [2:0] v_2599_0;
  wire [2:0] v_2600_0;
  reg [2:0] v_2601_0 = 3'h0;
  wire [0:0] v_2602_0;
  wire [0:0] v_2603_0;
  wire [0:0] v_2604_0;
  wire [2:0] v_2605_0;
  wire [2:0] v_2606_0;
  wire [2:0] v_2607_0;
  reg [2:0] v_2608_0 = 3'h0;
  wire [0:0] v_2609_0;
  wire [0:0] v_2610_0;
  wire [0:0] v_2611_0;
  wire [2:0] v_2612_0;
  wire [2:0] v_2613_0;
  wire [2:0] v_2614_0;
  reg [2:0] v_2615_0 = 3'h0;
  wire [0:0] v_2616_0;
  wire [0:0] v_2617_0;
  wire [0:0] v_2618_0;
  wire [2:0] v_2619_0;
  wire [2:0] v_2620_0;
  wire [2:0] v_2621_0;
  reg [2:0] v_2622_0 = 3'h0;
  wire [0:0] v_2623_0;
  wire [0:0] v_2624_0;
  wire [0:0] v_2625_0;
  wire [2:0] v_2626_0;
  wire [2:0] v_2627_0;
  wire [2:0] v_2628_0;
  reg [2:0] v_2629_0 = 3'h0;
  wire [0:0] v_2630_0;
  wire [0:0] v_2631_0;
  wire [0:0] v_2632_0;
  wire [2:0] v_2633_0;
  wire [2:0] v_2634_0;
  wire [2:0] v_2635_0;
  reg [2:0] v_2636_0 = 3'h0;
  wire [0:0] v_2637_0;
  wire [0:0] v_2638_0;
  wire [0:0] v_2639_0;
  wire [2:0] v_2640_0;
  wire [2:0] v_2641_0;
  wire [2:0] v_2642_0;
  reg [2:0] v_2643_0 = 3'h0;
  wire [0:0] v_2644_0;
  wire [0:0] v_2645_0;
  wire [0:0] v_2646_0;
  wire [2:0] v_2647_0;
  wire [2:0] v_2648_0;
  wire [2:0] v_2649_0;
  reg [2:0] v_2650_0 = 3'h0;
  wire [0:0] v_2651_0;
  wire [0:0] v_2652_0;
  wire [0:0] v_2653_0;
  wire [2:0] v_2654_0;
  wire [2:0] v_2655_0;
  wire [2:0] v_2656_0;
  reg [2:0] v_2657_0 = 3'h0;
  wire [0:0] v_2658_0;
  wire [0:0] v_2659_0;
  wire [0:0] v_2660_0;
  wire [2:0] v_2661_0;
  wire [2:0] v_2662_0;
  wire [2:0] v_2663_0;
  reg [2:0] v_2664_0 = 3'h0;
  wire [0:0] v_2665_0;
  wire [0:0] v_2666_0;
  wire [0:0] v_2667_0;
  wire [2:0] v_2668_0;
  wire [2:0] v_2669_0;
  wire [2:0] v_2670_0;
  reg [2:0] v_2671_0 = 3'h0;
  wire [0:0] v_2672_0;
  wire [0:0] v_2673_0;
  wire [0:0] v_2674_0;
  wire [2:0] v_2675_0;
  wire [2:0] v_2676_0;
  wire [2:0] v_2677_0;
  reg [2:0] v_2678_0 = 3'h0;
  wire [0:0] v_2679_0;
  wire [0:0] v_2680_0;
  wire [0:0] v_2681_0;
  wire [2:0] v_2682_0;
  wire [2:0] v_2683_0;
  wire [2:0] v_2684_0;
  reg [2:0] v_2685_0 = 3'h0;
  wire [0:0] v_2686_0;
  wire [0:0] v_2687_0;
  wire [0:0] v_2688_0;
  wire [2:0] v_2689_0;
  wire [2:0] v_2690_0;
  wire [2:0] v_2691_0;
  reg [2:0] v_2692_0 = 3'h0;
  wire [0:0] v_2693_0;
  wire [0:0] v_2694_0;
  wire [0:0] v_2695_0;
  wire [2:0] v_2696_0;
  wire [2:0] v_2697_0;
  wire [2:0] v_2698_0;
  reg [2:0] v_2699_0 = 3'h0;
  wire [0:0] v_2700_0;
  wire [0:0] v_2701_0;
  wire [0:0] v_2702_0;
  wire [2:0] v_2703_0;
  wire [2:0] v_2704_0;
  wire [2:0] v_2705_0;
  reg [2:0] v_2706_0 = 3'h0;
  wire [0:0] v_2707_0;
  wire [0:0] v_2708_0;
  wire [0:0] v_2709_0;
  wire [2:0] v_2710_0;
  wire [2:0] v_2711_0;
  wire [2:0] v_2712_0;
  reg [2:0] v_2713_0 = 3'h0;
  wire [0:0] v_2714_0;
  wire [0:0] v_2715_0;
  wire [0:0] v_2716_0;
  wire [2:0] v_2717_0;
  wire [2:0] v_2718_0;
  wire [2:0] v_2719_0;
  reg [2:0] v_2720_0 = 3'h0;
  wire [0:0] v_2721_0;
  wire [0:0] v_2722_0;
  wire [0:0] v_2723_0;
  wire [2:0] v_2724_0;
  wire [2:0] v_2725_0;
  wire [2:0] v_2726_0;
  reg [2:0] v_2727_0 = 3'h0;
  wire [0:0] v_2728_0;
  wire [0:0] v_2729_0;
  wire [0:0] v_2730_0;
  wire [2:0] v_2731_0;
  wire [2:0] v_2732_0;
  wire [2:0] v_2733_0;
  reg [2:0] v_2734_0 = 3'h0;
  wire [0:0] v_2735_0;
  wire [0:0] v_2736_0;
  wire [0:0] v_2737_0;
  wire [2:0] v_2738_0;
  wire [2:0] v_2739_0;
  wire [2:0] v_2740_0;
  reg [2:0] v_2741_0 = 3'h0;
  wire [0:0] v_2742_0;
  wire [0:0] v_2743_0;
  wire [0:0] v_2744_0;
  wire [2:0] v_2745_0;
  wire [2:0] v_2746_0;
  wire [2:0] v_2747_0;
  reg [2:0] v_2748_0 = 3'h0;
  wire [0:0] v_2749_0;
  wire [0:0] v_2750_0;
  wire [0:0] v_2751_0;
  wire [2:0] v_2752_0;
  wire [2:0] v_2753_0;
  wire [2:0] v_2754_0;
  reg [2:0] v_2755_0 = 3'h0;
  wire [0:0] v_2756_0;
  wire [0:0] v_2757_0;
  wire [0:0] v_2758_0;
  wire [2:0] v_2759_0;
  wire [2:0] v_2760_0;
  wire [2:0] v_2761_0;
  reg [2:0] v_2762_0 = 3'h0;
  wire [0:0] v_2763_0;
  wire [0:0] v_2764_0;
  wire [0:0] v_2765_0;
  wire [2:0] v_2766_0;
  wire [2:0] v_2767_0;
  wire [2:0] v_2768_0;
  reg [2:0] v_2769_0 = 3'h0;
  wire [0:0] v_2770_0;
  wire [0:0] v_2771_0;
  wire [0:0] v_2772_0;
  wire [2:0] v_2773_0;
  wire [2:0] v_2774_0;
  wire [2:0] v_2775_0;
  reg [2:0] v_2776_0 = 3'h0;
  wire [0:0] v_2777_0;
  wire [0:0] v_2778_0;
  wire [0:0] v_2779_0;
  wire [2:0] v_2780_0;
  wire [2:0] v_2781_0;
  wire [2:0] v_2782_0;
  reg [2:0] v_2783_0 = 3'h0;
  wire [0:0] v_2784_0;
  wire [0:0] v_2785_0;
  wire [0:0] v_2786_0;
  wire [2:0] v_2787_0;
  wire [2:0] v_2788_0;
  wire [2:0] v_2789_0;
  reg [2:0] v_2790_0 = 3'h0;
  wire [0:0] v_2791_0;
  wire [0:0] v_2792_0;
  wire [0:0] v_2793_0;
  wire [2:0] v_2794_0;
  wire [2:0] v_2795_0;
  wire [2:0] v_2796_0;
  reg [2:0] v_2797_0 = 3'h0;
  wire [0:0] v_2798_0;
  wire [0:0] v_2799_0;
  wire [0:0] v_2800_0;
  wire [2:0] v_2801_0;
  wire [2:0] v_2802_0;
  wire [2:0] v_2803_0;
  reg [2:0] v_2804_0 = 3'h0;
  wire [0:0] v_2805_0;
  wire [0:0] v_2806_0;
  wire [0:0] v_2807_0;
  wire [2:0] v_2808_0;
  wire [2:0] v_2809_0;
  wire [2:0] v_2810_0;
  reg [2:0] v_2811_0 = 3'h0;
  wire [0:0] v_2812_0;
  wire [0:0] v_2813_0;
  wire [0:0] v_2814_0;
  wire [2:0] v_2815_0;
  wire [2:0] v_2816_0;
  wire [2:0] v_2817_0;
  reg [2:0] v_2818_0 = 3'h0;
  wire [0:0] v_2819_0;
  wire [0:0] v_2820_0;
  wire [0:0] v_2821_0;
  wire [2:0] v_2822_0;
  wire [2:0] v_2823_0;
  wire [2:0] v_2824_0;
  reg [2:0] v_2825_0 = 3'h0;
  wire [0:0] v_2826_0;
  wire [0:0] v_2827_0;
  wire [0:0] v_2828_0;
  wire [2:0] v_2829_0;
  wire [2:0] v_2830_0;
  wire [2:0] v_2831_0;
  reg [2:0] v_2832_0 = 3'h0;
  wire [0:0] v_2833_0;
  wire [0:0] v_2834_0;
  wire [0:0] v_2835_0;
  wire [2:0] v_2836_0;
  wire [2:0] v_2837_0;
  wire [2:0] v_2838_0;
  reg [2:0] v_2839_0 = 3'h0;
  wire [0:0] v_2840_0;
  wire [0:0] v_2841_0;
  wire [0:0] v_2842_0;
  wire [2:0] v_2843_0;
  wire [2:0] v_2844_0;
  wire [2:0] v_2845_0;
  reg [2:0] v_2846_0 = 3'h0;
  wire [0:0] v_2847_0;
  wire [0:0] v_2848_0;
  wire [0:0] v_2849_0;
  wire [2:0] v_2850_0;
  wire [2:0] v_2851_0;
  wire [2:0] v_2852_0;
  reg [2:0] v_2853_0 = 3'h0;
  wire [0:0] v_2854_0;
  wire [0:0] v_2855_0;
  wire [0:0] v_2856_0;
  wire [2:0] v_2857_0;
  wire [2:0] v_2858_0;
  wire [2:0] v_2859_0;
  reg [2:0] v_2860_0 = 3'h0;
  wire [0:0] v_2861_0;
  wire [0:0] v_2862_0;
  wire [0:0] v_2863_0;
  wire [2:0] v_2864_0;
  wire [2:0] v_2865_0;
  wire [2:0] v_2866_0;
  reg [2:0] v_2867_0 = 3'h0;
  wire [0:0] v_2868_0;
  wire [0:0] v_2869_0;
  wire [0:0] v_2870_0;
  wire [2:0] v_2871_0;
  wire [2:0] v_2872_0;
  wire [2:0] v_2873_0;
  reg [2:0] v_2874_0 = 3'h0;
  wire [0:0] v_2875_0;
  wire [0:0] v_2876_0;
  wire [0:0] v_2877_0;
  wire [2:0] v_2878_0;
  wire [2:0] v_2879_0;
  wire [2:0] v_2880_0;
  reg [2:0] v_2881_0 = 3'h0;
  wire [0:0] v_2882_0;
  wire [0:0] v_2883_0;
  wire [0:0] v_2884_0;
  wire [2:0] v_2885_0;
  wire [2:0] v_2886_0;
  wire [2:0] v_2887_0;
  reg [2:0] v_2888_0 = 3'h0;
  wire [0:0] v_2889_0;
  wire [0:0] v_2890_0;
  wire [0:0] v_2891_0;
  wire [2:0] v_2892_0;
  wire [2:0] v_2893_0;
  wire [2:0] v_2894_0;
  reg [2:0] v_2895_0 = 3'h0;
  wire [0:0] v_2896_0;
  wire [0:0] v_2897_0;
  wire [0:0] v_2898_0;
  wire [2:0] v_2899_0;
  wire [2:0] v_2900_0;
  wire [2:0] v_2901_0;
  reg [2:0] v_2902_0 = 3'h0;
  wire [0:0] v_2903_0;
  wire [0:0] v_2904_0;
  wire [0:0] v_2905_0;
  wire [2:0] v_2906_0;
  wire [2:0] v_2907_0;
  wire [2:0] v_2908_0;
  reg [2:0] v_2909_0 = 3'h0;
  wire [0:0] v_2910_0;
  wire [0:0] v_2911_0;
  wire [0:0] v_2912_0;
  wire [2:0] v_2913_0;
  wire [2:0] v_2914_0;
  wire [2:0] v_2915_0;
  reg [2:0] v_2916_0 = 3'h0;
  wire [0:0] v_2917_0;
  wire [0:0] v_2918_0;
  wire [0:0] v_2919_0;
  wire [2:0] v_2920_0;
  wire [2:0] v_2921_0;
  wire [2:0] v_2922_0;
  reg [2:0] v_2923_0 = 3'h0;
  wire [0:0] v_2924_0;
  wire [0:0] v_2925_0;
  wire [0:0] v_2926_0;
  wire [2:0] v_2927_0;
  wire [2:0] v_2928_0;
  wire [2:0] v_2929_0;
  reg [2:0] v_2930_0 = 3'h0;
  wire [0:0] v_2931_0;
  wire [0:0] v_2932_0;
  wire [0:0] v_2933_0;
  wire [2:0] v_2934_0;
  wire [2:0] v_2935_0;
  wire [2:0] v_2936_0;
  reg [2:0] v_2937_0 = 3'h0;
  wire [0:0] v_2938_0;
  wire [0:0] v_2939_0;
  wire [0:0] v_2940_0;
  wire [2:0] v_2941_0;
  wire [2:0] v_2942_0;
  wire [2:0] v_2943_0;
  reg [2:0] v_2944_0 = 3'h0;
  wire [0:0] v_2945_0;
  wire [0:0] v_2946_0;
  wire [0:0] v_2947_0;
  wire [2:0] v_2948_0;
  wire [2:0] v_2949_0;
  wire [2:0] v_2950_0;
  reg [2:0] v_2951_0 = 3'h0;
  wire [0:0] v_2952_0;
  wire [0:0] v_2953_0;
  wire [0:0] v_2954_0;
  wire [2:0] v_2955_0;
  wire [2:0] v_2956_0;
  wire [2:0] v_2957_0;
  reg [2:0] v_2958_0 = 3'h0;
  wire [0:0] v_2959_0;
  wire [0:0] v_2960_0;
  wire [0:0] v_2961_0;
  wire [2:0] v_2962_0;
  wire [2:0] v_2963_0;
  wire [2:0] v_2964_0;
  reg [2:0] v_2965_0 = 3'h0;
  wire [0:0] v_2966_0;
  wire [0:0] v_2967_0;
  wire [0:0] v_2968_0;
  wire [2:0] v_2969_0;
  wire [2:0] v_2970_0;
  wire [2:0] v_2971_0;
  reg [2:0] v_2972_0 = 3'h0;
  wire [0:0] v_2973_0;
  wire [0:0] v_2974_0;
  wire [0:0] v_2975_0;
  wire [2:0] v_2976_0;
  wire [2:0] v_2977_0;
  wire [2:0] v_2978_0;
  reg [2:0] v_2979_0 = 3'h0;
  wire [0:0] v_2980_0;
  wire [0:0] v_2981_0;
  wire [0:0] v_2982_0;
  wire [2:0] v_2983_0;
  wire [2:0] v_2984_0;
  wire [2:0] v_2985_0;
  reg [2:0] v_2986_0 = 3'h0;
  wire [0:0] v_2987_0;
  wire [0:0] v_2988_0;
  wire [0:0] v_2989_0;
  wire [2:0] v_2990_0;
  wire [2:0] v_2991_0;
  wire [2:0] v_2992_0;
  reg [2:0] v_2993_0 = 3'h0;
  wire [0:0] v_2994_0;
  wire [0:0] v_2995_0;
  wire [0:0] v_2996_0;
  wire [2:0] v_2997_0;
  wire [2:0] v_2998_0;
  wire [2:0] v_2999_0;
  reg [2:0] v_3000_0 = 3'h0;
  wire [0:0] v_3001_0;
  wire [0:0] v_3002_0;
  wire [0:0] v_3003_0;
  wire [2:0] v_3004_0;
  wire [2:0] v_3005_0;
  wire [2:0] v_3006_0;
  reg [2:0] v_3007_0 = 3'h0;
  wire [0:0] v_3008_0;
  wire [0:0] v_3009_0;
  wire [0:0] v_3010_0;
  wire [2:0] v_3011_0;
  wire [2:0] v_3012_0;
  wire [2:0] v_3013_0;
  reg [2:0] v_3014_0 = 3'h0;
  wire [0:0] v_3015_0;
  wire [0:0] v_3016_0;
  wire [0:0] v_3017_0;
  wire [2:0] v_3018_0;
  wire [2:0] v_3019_0;
  wire [2:0] v_3020_0;
  reg [2:0] v_3021_0 = 3'h0;
  wire [0:0] v_3022_0;
  wire [0:0] v_3023_0;
  wire [0:0] v_3024_0;
  wire [2:0] v_3025_0;
  wire [2:0] v_3026_0;
  wire [2:0] v_3027_0;
  reg [2:0] v_3028_0 = 3'h0;
  wire [0:0] v_3029_0;
  wire [0:0] v_3030_0;
  wire [0:0] v_3031_0;
  wire [2:0] v_3032_0;
  wire [2:0] v_3033_0;
  wire [2:0] v_3034_0;
  reg [2:0] v_3035_0 = 3'h0;
  wire [0:0] v_3036_0;
  wire [0:0] v_3037_0;
  wire [0:0] v_3038_0;
  wire [2:0] v_3039_0;
  wire [2:0] v_3040_0;
  wire [2:0] v_3041_0;
  reg [2:0] v_3042_0 = 3'h0;
  wire [0:0] v_3043_0;
  wire [0:0] v_3044_0;
  wire [0:0] v_3045_0;
  wire [2:0] v_3046_0;
  wire [2:0] v_3047_0;
  wire [2:0] v_3048_0;
  reg [2:0] v_3049_0 = 3'h0;
  wire [0:0] v_3050_0;
  wire [0:0] v_3051_0;
  wire [0:0] v_3052_0;
  wire [2:0] v_3053_0;
  wire [2:0] v_3054_0;
  wire [2:0] v_3055_0;
  reg [2:0] v_3056_0 = 3'h0;
  wire [0:0] v_3057_0;
  wire [0:0] v_3058_0;
  wire [0:0] v_3059_0;
  wire [2:0] v_3060_0;
  wire [2:0] v_3061_0;
  wire [2:0] v_3062_0;
  reg [2:0] v_3063_0 = 3'h0;
  wire [0:0] v_3064_0;
  wire [0:0] v_3065_0;
  wire [0:0] v_3066_0;
  wire [2:0] v_3067_0;
  wire [2:0] v_3068_0;
  wire [2:0] v_3069_0;
  reg [2:0] v_3070_0 = 3'h0;
  wire [0:0] v_3071_0;
  wire [0:0] v_3072_0;
  wire [0:0] v_3073_0;
  wire [2:0] v_3074_0;
  wire [2:0] v_3075_0;
  wire [2:0] v_3076_0;
  reg [2:0] v_3077_0 = 3'h0;
  wire [0:0] v_3078_0;
  wire [0:0] v_3079_0;
  wire [0:0] v_3080_0;
  wire [2:0] v_3081_0;
  wire [2:0] v_3082_0;
  wire [2:0] v_3083_0;
  reg [2:0] v_3084_0 = 3'h0;
  wire [0:0] v_3085_0;
  wire [0:0] v_3086_0;
  wire [0:0] v_3087_0;
  wire [2:0] v_3088_0;
  wire [2:0] v_3089_0;
  wire [2:0] v_3090_0;
  reg [2:0] v_3091_0 = 3'h0;
  wire [0:0] v_3092_0;
  wire [0:0] v_3093_0;
  wire [0:0] v_3094_0;
  wire [2:0] v_3095_0;
  wire [2:0] v_3096_0;
  wire [2:0] v_3097_0;
  reg [2:0] v_3098_0 = 3'h0;
  wire [0:0] v_3099_0;
  wire [0:0] v_3100_0;
  wire [0:0] v_3101_0;
  wire [2:0] v_3102_0;
  wire [2:0] v_3103_0;
  wire [2:0] v_3104_0;
  reg [2:0] v_3105_0 = 3'h0;
  wire [0:0] v_3106_0;
  wire [0:0] v_3107_0;
  wire [0:0] v_3108_0;
  wire [2:0] v_3109_0;
  wire [2:0] v_3110_0;
  wire [2:0] v_3111_0;
  reg [2:0] v_3112_0 = 3'h0;
  wire [0:0] v_3113_0;
  wire [0:0] v_3114_0;
  wire [0:0] v_3115_0;
  wire [2:0] v_3116_0;
  wire [2:0] v_3117_0;
  wire [2:0] v_3118_0;
  reg [2:0] v_3119_0 = 3'h0;
  wire [0:0] v_3120_0;
  wire [0:0] v_3121_0;
  wire [0:0] v_3122_0;
  wire [2:0] v_3123_0;
  wire [2:0] v_3124_0;
  wire [2:0] v_3125_0;
  reg [2:0] v_3126_0 = 3'h0;
  wire [0:0] v_3127_0;
  wire [0:0] v_3128_0;
  wire [0:0] v_3129_0;
  wire [2:0] v_3130_0;
  wire [2:0] v_3131_0;
  wire [2:0] v_3132_0;
  reg [2:0] v_3133_0 = 3'h0;
  wire [0:0] v_3134_0;
  wire [0:0] v_3135_0;
  wire [0:0] v_3136_0;
  wire [2:0] v_3137_0;
  wire [2:0] v_3138_0;
  wire [2:0] v_3139_0;
  reg [2:0] v_3140_0 = 3'h0;
  wire [0:0] v_3141_0;
  wire [0:0] v_3142_0;
  wire [0:0] v_3143_0;
  wire [2:0] v_3144_0;
  wire [2:0] v_3145_0;
  wire [2:0] v_3146_0;
  reg [2:0] v_3147_0 = 3'h0;
  wire [0:0] v_3148_0;
  wire [0:0] v_3149_0;
  wire [0:0] v_3150_0;
  wire [2:0] v_3151_0;
  wire [2:0] v_3152_0;
  wire [2:0] v_3153_0;
  reg [2:0] v_3154_0 = 3'h0;
  wire [0:0] v_3155_0;
  wire [0:0] v_3156_0;
  wire [0:0] v_3157_0;
  wire [2:0] v_3158_0;
  wire [2:0] v_3159_0;
  wire [2:0] v_3160_0;
  reg [2:0] v_3161_0 = 3'h0;
  wire [0:0] v_3162_0;
  wire [0:0] v_3163_0;
  wire [0:0] v_3164_0;
  wire [2:0] v_3165_0;
  wire [2:0] v_3166_0;
  wire [2:0] v_3167_0;
  reg [2:0] v_3168_0 = 3'h0;
  wire [0:0] v_3169_0;
  wire [0:0] v_3170_0;
  wire [0:0] v_3171_0;
  wire [2:0] v_3172_0;
  wire [2:0] v_3173_0;
  wire [2:0] v_3174_0;
  reg [2:0] v_3175_0 = 3'h0;
  wire [0:0] v_3176_0;
  wire [0:0] v_3177_0;
  wire [0:0] v_3178_0;
  wire [2:0] v_3179_0;
  wire [2:0] v_3180_0;
  wire [2:0] v_3181_0;
  reg [2:0] v_3182_0 = 3'h0;
  wire [0:0] v_3183_0;
  wire [0:0] v_3184_0;
  wire [0:0] v_3185_0;
  wire [2:0] v_3186_0;
  wire [2:0] v_3187_0;
  wire [2:0] v_3188_0;
  reg [2:0] v_3189_0 = 3'h0;
  wire [0:0] v_3190_0;
  wire [0:0] v_3191_0;
  wire [0:0] v_3192_0;
  wire [2:0] v_3193_0;
  wire [2:0] v_3194_0;
  wire [2:0] v_3195_0;
  reg [2:0] v_3196_0 = 3'h0;
  wire [0:0] v_3197_0;
  wire [0:0] v_3198_0;
  wire [0:0] v_3199_0;
  wire [2:0] v_3200_0;
  wire [2:0] v_3201_0;
  wire [2:0] v_3202_0;
  reg [2:0] v_3203_0 = 3'h0;
  wire [0:0] v_3204_0;
  wire [0:0] v_3205_0;
  wire [0:0] v_3206_0;
  wire [2:0] v_3207_0;
  wire [2:0] v_3208_0;
  wire [2:0] v_3209_0;
  reg [2:0] v_3210_0 = 3'h0;
  wire [0:0] v_3211_0;
  wire [0:0] v_3212_0;
  wire [0:0] v_3213_0;
  wire [2:0] v_3214_0;
  wire [2:0] v_3215_0;
  wire [2:0] v_3216_0;
  reg [2:0] v_3217_0 = 3'h0;
  wire [0:0] v_3218_0;
  wire [0:0] v_3219_0;
  wire [0:0] v_3220_0;
  wire [2:0] v_3221_0;
  wire [2:0] v_3222_0;
  wire [2:0] v_3223_0;
  reg [2:0] v_3224_0 = 3'h0;
  wire [0:0] v_3225_0;
  wire [0:0] v_3226_0;
  wire [0:0] v_3227_0;
  wire [2:0] v_3228_0;
  wire [2:0] v_3229_0;
  wire [2:0] v_3230_0;
  reg [2:0] v_3231_0 = 3'h0;
  wire [0:0] v_3232_0;
  wire [0:0] v_3233_0;
  wire [0:0] v_3234_0;
  wire [2:0] v_3235_0;
  wire [2:0] v_3236_0;
  wire [2:0] v_3237_0;
  reg [2:0] v_3238_0 = 3'h0;
  wire [0:0] v_3239_0;
  wire [0:0] v_3240_0;
  wire [0:0] v_3241_0;
  wire [2:0] v_3242_0;
  wire [2:0] v_3243_0;
  wire [2:0] v_3244_0;
  reg [2:0] v_3245_0 = 3'h0;
  wire [0:0] v_3246_0;
  wire [0:0] v_3247_0;
  wire [0:0] v_3248_0;
  wire [2:0] v_3249_0;
  wire [2:0] v_3250_0;
  wire [2:0] v_3251_0;
  reg [2:0] v_3252_0 = 3'h0;
  wire [0:0] v_3253_0;
  wire [0:0] v_3254_0;
  wire [0:0] v_3255_0;
  wire [2:0] v_3256_0;
  wire [2:0] v_3257_0;
  wire [2:0] v_3258_0;
  reg [2:0] v_3259_0 = 3'h0;
  wire [0:0] v_3260_0;
  wire [0:0] v_3261_0;
  wire [0:0] v_3262_0;
  wire [2:0] v_3263_0;
  wire [2:0] v_3264_0;
  wire [2:0] v_3265_0;
  reg [2:0] v_3266_0 = 3'h0;
  wire [0:0] v_3267_0;
  wire [0:0] v_3268_0;
  wire [0:0] v_3269_0;
  wire [2:0] v_3270_0;
  wire [2:0] v_3271_0;
  wire [2:0] v_3272_0;
  reg [2:0] v_3273_0 = 3'h0;
  wire [0:0] v_3274_0;
  wire [0:0] v_3275_0;
  wire [0:0] v_3276_0;
  wire [2:0] v_3277_0;
  wire [2:0] v_3278_0;
  wire [2:0] v_3279_0;
  reg [2:0] v_3280_0 = 3'h0;
  wire [0:0] v_3281_0;
  wire [0:0] v_3282_0;
  wire [0:0] v_3283_0;
  wire [2:0] v_3284_0;
  wire [2:0] v_3285_0;
  wire [2:0] v_3286_0;
  reg [2:0] v_3287_0 = 3'h0;
  wire [0:0] v_3288_0;
  wire [0:0] v_3289_0;
  wire [0:0] v_3290_0;
  wire [2:0] v_3291_0;
  wire [2:0] v_3292_0;
  wire [2:0] v_3293_0;
  reg [2:0] v_3294_0 = 3'h0;
  wire [0:0] v_3295_0;
  wire [0:0] v_3296_0;
  wire [0:0] v_3297_0;
  wire [2:0] v_3298_0;
  wire [2:0] v_3299_0;
  wire [2:0] v_3300_0;
  reg [2:0] v_3301_0 = 3'h0;
  wire [0:0] v_3302_0;
  wire [0:0] v_3303_0;
  wire [0:0] v_3304_0;
  wire [2:0] v_3305_0;
  wire [2:0] v_3306_0;
  wire [2:0] v_3307_0;
  reg [2:0] v_3308_0 = 3'h0;
  wire [0:0] v_3309_0;
  wire [0:0] v_3310_0;
  wire [0:0] v_3311_0;
  wire [2:0] v_3312_0;
  wire [2:0] v_3313_0;
  wire [2:0] v_3314_0;
  reg [2:0] v_3315_0 = 3'h0;
  wire [0:0] v_3316_0;
  wire [0:0] v_3317_0;
  wire [0:0] v_3318_0;
  wire [2:0] v_3319_0;
  wire [2:0] v_3320_0;
  wire [2:0] v_3321_0;
  reg [2:0] v_3322_0 = 3'h0;
  wire [0:0] v_3323_0;
  wire [0:0] v_3324_0;
  wire [0:0] v_3325_0;
  wire [2:0] v_3326_0;
  wire [2:0] v_3327_0;
  wire [2:0] v_3328_0;
  reg [2:0] v_3329_0 = 3'h0;
  wire [0:0] v_3330_0;
  wire [0:0] v_3331_0;
  wire [0:0] v_3332_0;
  wire [2:0] v_3333_0;
  wire [2:0] v_3334_0;
  wire [2:0] v_3335_0;
  reg [2:0] v_3336_0 = 3'h0;
  wire [0:0] v_3337_0;
  wire [0:0] v_3338_0;
  wire [0:0] v_3339_0;
  wire [2:0] v_3340_0;
  wire [2:0] v_3341_0;
  wire [2:0] v_3342_0;
  reg [2:0] v_3343_0 = 3'h0;
  wire [0:0] v_3344_0;
  wire [0:0] v_3345_0;
  wire [0:0] v_3346_0;
  wire [2:0] v_3347_0;
  wire [2:0] v_3348_0;
  wire [2:0] v_3349_0;
  reg [2:0] v_3350_0 = 3'h0;
  wire [0:0] v_3351_0;
  wire [0:0] v_3352_0;
  wire [0:0] v_3353_0;
  wire [2:0] v_3354_0;
  wire [2:0] v_3355_0;
  wire [2:0] v_3356_0;
  reg [2:0] v_3357_0 = 3'h0;
  wire [0:0] v_3358_0;
  wire [0:0] v_3359_0;
  wire [0:0] v_3360_0;
  wire [2:0] v_3361_0;
  wire [2:0] v_3362_0;
  wire [2:0] v_3363_0;
  reg [2:0] v_3364_0 = 3'h0;
  wire [0:0] v_3365_0;
  wire [0:0] v_3366_0;
  wire [0:0] v_3367_0;
  wire [2:0] v_3368_0;
  wire [2:0] v_3369_0;
  wire [2:0] v_3370_0;
  reg [2:0] v_3371_0 = 3'h0;
  wire [0:0] v_3372_0;
  wire [0:0] v_3373_0;
  wire [0:0] v_3374_0;
  wire [2:0] v_3375_0;
  wire [2:0] v_3376_0;
  wire [2:0] v_3377_0;
  reg [2:0] v_3378_0 = 3'h0;
  wire [0:0] v_3379_0;
  wire [0:0] v_3380_0;
  wire [0:0] v_3381_0;
  wire [2:0] v_3382_0;
  wire [2:0] v_3383_0;
  wire [2:0] v_3384_0;
  reg [2:0] v_3385_0 = 3'h0;
  wire [0:0] v_3386_0;
  wire [0:0] v_3387_0;
  wire [0:0] v_3388_0;
  wire [2:0] v_3389_0;
  wire [2:0] v_3390_0;
  wire [2:0] v_3391_0;
  reg [2:0] v_3392_0 = 3'h0;
  wire [0:0] v_3393_0;
  wire [0:0] v_3394_0;
  wire [0:0] v_3395_0;
  wire [2:0] v_3396_0;
  wire [2:0] v_3397_0;
  wire [2:0] v_3398_0;
  reg [2:0] v_3399_0 = 3'h0;
  wire [0:0] v_3400_0;
  wire [0:0] v_3401_0;
  wire [0:0] v_3402_0;
  wire [2:0] v_3403_0;
  wire [2:0] v_3404_0;
  wire [2:0] v_3405_0;
  reg [2:0] v_3406_0 = 3'h0;
  wire [0:0] v_3407_0;
  wire [0:0] v_3408_0;
  wire [0:0] v_3409_0;
  wire [2:0] v_3410_0;
  wire [2:0] v_3411_0;
  wire [2:0] v_3412_0;
  reg [2:0] v_3413_0 = 3'h0;
  wire [0:0] v_3414_0;
  wire [0:0] v_3415_0;
  wire [0:0] v_3416_0;
  wire [2:0] v_3417_0;
  wire [2:0] v_3418_0;
  wire [2:0] v_3419_0;
  reg [2:0] v_3420_0 = 3'h0;
  wire [0:0] v_3421_0;
  wire [0:0] v_3422_0;
  wire [0:0] v_3423_0;
  wire [2:0] v_3424_0;
  wire [2:0] v_3425_0;
  wire [2:0] v_3426_0;
  reg [2:0] v_3427_0 = 3'h0;
  wire [0:0] v_3428_0;
  wire [0:0] v_3429_0;
  wire [0:0] v_3430_0;
  wire [2:0] v_3431_0;
  wire [2:0] v_3432_0;
  wire [2:0] v_3433_0;
  reg [2:0] v_3434_0 = 3'h0;
  wire [0:0] v_3435_0;
  wire [0:0] v_3436_0;
  wire [0:0] v_3437_0;
  wire [2:0] v_3438_0;
  wire [2:0] v_3439_0;
  wire [2:0] v_3440_0;
  reg [2:0] v_3441_0 = 3'h0;
  wire [0:0] v_3442_0;
  wire [0:0] v_3443_0;
  wire [0:0] v_3444_0;
  wire [2:0] v_3445_0;
  wire [2:0] v_3446_0;
  wire [2:0] v_3447_0;
  reg [2:0] v_3448_0 = 3'h0;
  wire [0:0] v_3449_0;
  wire [0:0] v_3450_0;
  wire [0:0] v_3451_0;
  wire [2:0] v_3452_0;
  wire [2:0] v_3453_0;
  wire [2:0] v_3454_0;
  reg [2:0] v_3455_0 = 3'h0;
  wire [0:0] v_3456_0;
  wire [0:0] v_3457_0;
  wire [0:0] v_3458_0;
  wire [2:0] v_3459_0;
  wire [2:0] v_3460_0;
  wire [2:0] v_3461_0;
  reg [2:0] v_3462_0 = 3'h0;
  wire [0:0] v_3463_0;
  wire [0:0] v_3464_0;
  wire [0:0] v_3465_0;
  wire [2:0] v_3466_0;
  wire [2:0] v_3467_0;
  wire [2:0] v_3468_0;
  reg [2:0] v_3469_0 = 3'h0;
  wire [0:0] v_3470_0;
  wire [0:0] v_3471_0;
  wire [0:0] v_3472_0;
  wire [2:0] v_3473_0;
  wire [2:0] v_3474_0;
  wire [2:0] v_3475_0;
  reg [2:0] v_3476_0 = 3'h0;
  wire [0:0] v_3477_0;
  wire [0:0] v_3478_0;
  wire [0:0] v_3479_0;
  wire [2:0] v_3480_0;
  wire [2:0] v_3481_0;
  wire [2:0] v_3482_0;
  reg [2:0] v_3483_0 = 3'h0;
  wire [0:0] v_3484_0;
  wire [0:0] v_3485_0;
  wire [0:0] v_3486_0;
  wire [2:0] v_3487_0;
  wire [2:0] v_3488_0;
  wire [2:0] v_3489_0;
  reg [2:0] v_3490_0 = 3'h0;
  wire [0:0] v_3491_0;
  wire [0:0] v_3492_0;
  wire [0:0] v_3493_0;
  wire [2:0] v_3494_0;
  wire [2:0] v_3495_0;
  wire [2:0] v_3496_0;
  reg [2:0] v_3497_0 = 3'h0;
  wire [0:0] v_3498_0;
  wire [0:0] v_3499_0;
  wire [0:0] v_3500_0;
  wire [2:0] v_3501_0;
  wire [2:0] v_3502_0;
  wire [2:0] v_3503_0;
  reg [2:0] v_3504_0 = 3'h0;
  wire [0:0] v_3505_0;
  wire [0:0] v_3506_0;
  wire [0:0] v_3507_0;
  wire [2:0] v_3508_0;
  wire [2:0] v_3509_0;
  wire [2:0] v_3510_0;
  reg [2:0] v_3511_0 = 3'h0;
  wire [0:0] v_3512_0;
  wire [0:0] v_3513_0;
  wire [0:0] v_3514_0;
  wire [2:0] v_3515_0;
  wire [2:0] v_3516_0;
  wire [2:0] v_3517_0;
  reg [2:0] v_3518_0 = 3'h0;
  wire [0:0] v_3519_0;
  wire [0:0] v_3520_0;
  wire [0:0] v_3521_0;
  wire [2:0] v_3522_0;
  wire [2:0] v_3523_0;
  wire [2:0] v_3524_0;
  reg [2:0] v_3525_0 = 3'h0;
  wire [0:0] v_3526_0;
  wire [0:0] v_3527_0;
  wire [0:0] v_3528_0;
  wire [2:0] v_3529_0;
  wire [2:0] v_3530_0;
  wire [2:0] v_3531_0;
  reg [2:0] v_3532_0 = 3'h0;
  wire [0:0] v_3533_0;
  wire [0:0] v_3534_0;
  wire [0:0] v_3535_0;
  wire [2:0] v_3536_0;
  wire [2:0] v_3537_0;
  wire [2:0] v_3538_0;
  reg [2:0] v_3539_0 = 3'h0;
  wire [0:0] v_3540_0;
  wire [0:0] v_3541_0;
  wire [0:0] v_3542_0;
  wire [2:0] v_3543_0;
  wire [2:0] v_3544_0;
  wire [2:0] v_3545_0;
  reg [2:0] v_3546_0 = 3'h0;
  wire [0:0] v_3547_0;
  wire [0:0] v_3548_0;
  wire [0:0] v_3549_0;
  wire [2:0] v_3550_0;
  wire [2:0] v_3551_0;
  wire [2:0] v_3552_0;
  reg [2:0] v_3553_0 = 3'h0;
  wire [0:0] v_3554_0;
  wire [0:0] v_3555_0;
  wire [0:0] v_3556_0;
  wire [2:0] v_3557_0;
  wire [2:0] v_3558_0;
  wire [2:0] v_3559_0;
  reg [2:0] v_3560_0 = 3'h0;
  wire [0:0] v_3561_0;
  wire [0:0] v_3562_0;
  wire [0:0] v_3563_0;
  wire [2:0] v_3564_0;
  wire [2:0] v_3565_0;
  wire [2:0] v_3566_0;
  reg [2:0] v_3567_0 = 3'h0;
  wire [0:0] v_3568_0;
  wire [0:0] v_3569_0;
  wire [0:0] v_3570_0;
  wire [2:0] v_3571_0;
  wire [2:0] v_3572_0;
  wire [2:0] v_3573_0;
  reg [2:0] v_3574_0 = 3'h0;
  wire [0:0] v_3575_0;
  wire [0:0] v_3576_0;
  wire [0:0] v_3577_0;
  wire [2:0] v_3578_0;
  wire [2:0] v_3579_0;
  wire [2:0] v_3580_0;
  reg [2:0] v_3581_0 = 3'h0;
  wire [0:0] v_3582_0;
  wire [0:0] v_3583_0;
  wire [0:0] v_3584_0;
  wire [2:0] v_3585_0;
  wire [2:0] v_3586_0;
  wire [2:0] v_3587_0;
  reg [2:0] v_3588_0 = 3'h0;
  wire [0:0] v_3589_0;
  wire [0:0] v_3590_0;
  wire [0:0] v_3591_0;
  wire [2:0] v_3592_0;
  wire [2:0] v_3593_0;
  wire [2:0] v_3594_0;
  reg [2:0] v_3595_0 = 3'h0;
  wire [0:0] v_3596_0;
  wire [0:0] v_3597_0;
  wire [0:0] v_3598_0;
  wire [2:0] v_3599_0;
  wire [2:0] v_3600_0;
  wire [2:0] v_3601_0;
  reg [2:0] v_3602_0 = 3'h0;
  wire [0:0] v_3603_0;
  wire [0:0] v_3604_0;
  wire [0:0] v_3605_0;
  wire [2:0] v_3606_0;
  wire [2:0] v_3607_0;
  wire [2:0] v_3608_0;
  reg [2:0] v_3609_0 = 3'h0;
  wire [0:0] v_3610_0;
  wire [0:0] v_3611_0;
  wire [0:0] v_3612_0;
  wire [2:0] v_3613_0;
  wire [2:0] v_3614_0;
  wire [2:0] v_3615_0;
  reg [2:0] v_3616_0 = 3'h0;
  wire [0:0] v_3617_0;
  wire [0:0] v_3618_0;
  wire [0:0] v_3619_0;
  wire [2:0] v_3620_0;
  wire [2:0] v_3621_0;
  wire [2:0] v_3622_0;
  reg [2:0] v_3623_0 = 3'h0;
  wire [0:0] v_3624_0;
  wire [0:0] v_3625_0;
  wire [0:0] v_3626_0;
  wire [2:0] v_3627_0;
  wire [2:0] v_3628_0;
  wire [2:0] v_3629_0;
  reg [2:0] v_3630_0 = 3'h0;
  wire [0:0] v_3631_0;
  wire [0:0] v_3632_0;
  wire [0:0] v_3633_0;
  wire [2:0] v_3634_0;
  wire [2:0] v_3635_0;
  wire [2:0] v_3636_0;
  reg [2:0] v_3637_0 = 3'h0;
  wire [0:0] v_3638_0;
  wire [0:0] v_3639_0;
  wire [0:0] v_3640_0;
  wire [2:0] v_3641_0;
  wire [2:0] v_3642_0;
  wire [2:0] v_3643_0;
  reg [2:0] v_3644_0 = 3'h0;
  wire [0:0] v_3645_0;
  wire [0:0] v_3646_0;
  wire [0:0] v_3647_0;
  wire [2:0] v_3648_0;
  wire [2:0] v_3649_0;
  wire [2:0] v_3650_0;
  reg [2:0] v_3651_0 = 3'h0;
  wire [0:0] v_3652_0;
  wire [0:0] v_3653_0;
  wire [0:0] v_3654_0;
  wire [2:0] v_3655_0;
  wire [2:0] v_3656_0;
  wire [2:0] v_3657_0;
  reg [2:0] v_3658_0 = 3'h0;
  wire [0:0] v_3659_0;
  wire [0:0] v_3660_0;
  wire [0:0] v_3661_0;
  wire [2:0] v_3662_0;
  wire [2:0] v_3663_0;
  wire [2:0] v_3664_0;
  reg [2:0] v_3665_0 = 3'h0;
  wire [0:0] v_3666_0;
  wire [0:0] v_3667_0;
  wire [0:0] v_3668_0;
  wire [2:0] v_3669_0;
  wire [2:0] v_3670_0;
  wire [2:0] v_3671_0;
  reg [2:0] v_3672_0 = 3'h0;
  wire [0:0] v_3673_0;
  wire [0:0] v_3674_0;
  wire [0:0] v_3675_0;
  wire [2:0] v_3676_0;
  wire [2:0] v_3677_0;
  wire [2:0] v_3678_0;
  reg [2:0] v_3679_0 = 3'h0;
  wire [0:0] v_3680_0;
  wire [0:0] v_3681_0;
  wire [0:0] v_3682_0;
  wire [2:0] v_3683_0;
  wire [2:0] v_3684_0;
  wire [2:0] v_3685_0;
  reg [2:0] v_3686_0 = 3'h0;
  wire [0:0] v_3687_0;
  wire [0:0] v_3688_0;
  wire [0:0] v_3689_0;
  wire [2:0] v_3690_0;
  wire [2:0] v_3691_0;
  wire [2:0] v_3692_0;
  reg [2:0] v_3693_0 = 3'h0;
  wire [0:0] v_3694_0;
  wire [0:0] v_3695_0;
  wire [0:0] v_3696_0;
  wire [2:0] v_3697_0;
  wire [2:0] v_3698_0;
  wire [2:0] v_3699_0;
  reg [2:0] v_3700_0 = 3'h0;
  wire [0:0] v_3701_0;
  wire [0:0] v_3702_0;
  wire [0:0] v_3703_0;
  wire [2:0] v_3704_0;
  wire [2:0] v_3705_0;
  wire [2:0] v_3706_0;
  reg [2:0] v_3707_0 = 3'h0;
  wire [0:0] v_3708_0;
  wire [0:0] v_3709_0;
  wire [0:0] v_3710_0;
  wire [2:0] v_3711_0;
  wire [2:0] v_3712_0;
  wire [2:0] v_3713_0;
  reg [2:0] v_3714_0 = 3'h0;
  wire [0:0] v_3715_0;
  wire [0:0] v_3716_0;
  wire [0:0] v_3717_0;
  wire [2:0] v_3718_0;
  wire [2:0] v_3719_0;
  wire [2:0] v_3720_0;
  reg [2:0] v_3721_0 = 3'h0;
  wire [0:0] v_3722_0;
  wire [0:0] v_3723_0;
  wire [0:0] v_3724_0;
  wire [2:0] v_3725_0;
  wire [2:0] v_3726_0;
  wire [2:0] v_3727_0;
  reg [2:0] v_3728_0 = 3'h0;
  wire [0:0] v_3729_0;
  wire [0:0] v_3730_0;
  wire [0:0] v_3731_0;
  wire [2:0] v_3732_0;
  wire [2:0] v_3733_0;
  wire [2:0] v_3734_0;
  reg [2:0] v_3735_0 = 3'h0;
  wire [0:0] v_3736_0;
  wire [0:0] v_3737_0;
  wire [0:0] v_3738_0;
  wire [2:0] v_3739_0;
  wire [2:0] v_3740_0;
  wire [2:0] v_3741_0;
  reg [2:0] v_3742_0 = 3'h0;
  wire [0:0] v_3743_0;
  wire [0:0] v_3744_0;
  wire [0:0] v_3745_0;
  wire [2:0] v_3746_0;
  wire [2:0] v_3747_0;
  wire [2:0] v_3748_0;
  reg [2:0] v_3749_0 = 3'h0;
  wire [0:0] v_3750_0;
  wire [0:0] v_3751_0;
  wire [0:0] v_3752_0;
  wire [2:0] v_3753_0;
  wire [2:0] v_3754_0;
  wire [2:0] v_3755_0;
  reg [2:0] v_3756_0 = 3'h0;
  wire [0:0] v_3757_0;
  wire [0:0] v_3758_0;
  wire [0:0] v_3759_0;
  wire [2:0] v_3760_0;
  wire [2:0] v_3761_0;
  wire [2:0] v_3762_0;
  reg [2:0] v_3763_0 = 3'h0;
  wire [0:0] v_3764_0;
  wire [0:0] v_3765_0;
  wire [0:0] v_3766_0;
  wire [2:0] v_3767_0;
  wire [2:0] v_3768_0;
  wire [2:0] v_3769_0;
  reg [2:0] v_3770_0 = 3'h0;
  wire [0:0] v_3771_0;
  wire [0:0] v_3772_0;
  wire [0:0] v_3773_0;
  wire [2:0] v_3774_0;
  wire [2:0] v_3775_0;
  wire [2:0] v_3776_0;
  reg [2:0] v_3777_0 = 3'h0;
  wire [0:0] v_3778_0;
  wire [0:0] v_3779_0;
  wire [0:0] v_3780_0;
  wire [2:0] v_3781_0;
  wire [2:0] v_3782_0;
  wire [2:0] v_3783_0;
  reg [2:0] v_3784_0 = 3'h0;
  wire [0:0] v_3785_0;
  wire [0:0] v_3786_0;
  wire [0:0] v_3787_0;
  wire [2:0] v_3788_0;
  wire [2:0] v_3789_0;
  wire [2:0] v_3790_0;
  reg [2:0] v_3791_0 = 3'h0;
  wire [0:0] v_3792_0;
  wire [0:0] v_3793_0;
  wire [0:0] v_3794_0;
  wire [2:0] v_3795_0;
  wire [2:0] v_3796_0;
  wire [2:0] v_3797_0;
  reg [2:0] v_3798_0 = 3'h0;
  wire [0:0] v_3799_0;
  wire [0:0] v_3800_0;
  wire [0:0] v_3801_0;
  wire [2:0] v_3802_0;
  wire [2:0] v_3803_0;
  wire [2:0] v_3804_0;
  reg [2:0] v_3805_0 = 3'h0;
  wire [0:0] v_3806_0;
  wire [0:0] v_3807_0;
  wire [0:0] v_3808_0;
  wire [2:0] v_3809_0;
  wire [2:0] v_3810_0;
  wire [2:0] v_3811_0;
  reg [2:0] v_3812_0 = 3'h0;
  wire [0:0] v_3813_0;
  wire [0:0] v_3814_0;
  wire [0:0] v_3815_0;
  wire [2:0] v_3816_0;
  wire [2:0] v_3817_0;
  wire [2:0] v_3818_0;
  reg [2:0] v_3819_0 = 3'h0;
  wire [0:0] v_3820_0;
  wire [0:0] v_3821_0;
  wire [0:0] v_3822_0;
  wire [2:0] v_3823_0;
  wire [2:0] v_3824_0;
  wire [2:0] v_3825_0;
  reg [2:0] v_3826_0 = 3'h0;
  wire [0:0] v_3827_0;
  wire [0:0] v_3828_0;
  wire [0:0] v_3829_0;
  wire [2:0] v_3830_0;
  wire [2:0] v_3831_0;
  wire [2:0] v_3832_0;
  reg [2:0] v_3833_0 = 3'h0;
  wire [0:0] v_3834_0;
  wire [0:0] v_3835_0;
  wire [0:0] v_3836_0;
  wire [2:0] v_3837_0;
  wire [2:0] v_3838_0;
  wire [2:0] v_3839_0;
  reg [2:0] v_3840_0 = 3'h0;
  wire [0:0] v_3841_0;
  wire [0:0] v_3842_0;
  wire [0:0] v_3843_0;
  wire [2:0] v_3844_0;
  wire [2:0] v_3845_0;
  wire [2:0] v_3846_0;
  reg [2:0] v_3847_0 = 3'h0;
  wire [0:0] v_3848_0;
  wire [0:0] v_3849_0;
  wire [0:0] v_3850_0;
  wire [2:0] v_3851_0;
  wire [2:0] v_3852_0;
  wire [2:0] v_3853_0;
  reg [2:0] v_3854_0 = 3'h0;
  wire [0:0] v_3855_0;
  wire [0:0] v_3856_0;
  wire [0:0] v_3857_0;
  wire [2:0] v_3858_0;
  wire [2:0] v_3859_0;
  wire [2:0] v_3860_0;
  reg [2:0] v_3861_0 = 3'h0;
  wire [0:0] v_3862_0;
  wire [0:0] v_3863_0;
  wire [0:0] v_3864_0;
  wire [2:0] v_3865_0;
  wire [2:0] v_3866_0;
  wire [2:0] v_3867_0;
  reg [2:0] v_3868_0 = 3'h0;
  wire [0:0] v_3869_0;
  wire [0:0] v_3870_0;
  wire [0:0] v_3871_0;
  wire [2:0] v_3872_0;
  wire [2:0] v_3873_0;
  wire [2:0] v_3874_0;
  reg [2:0] v_3875_0 = 3'h0;
  wire [0:0] v_3876_0;
  wire [0:0] v_3877_0;
  wire [0:0] v_3878_0;
  wire [2:0] v_3879_0;
  wire [2:0] v_3880_0;
  wire [2:0] v_3881_0;
  reg [2:0] v_3882_0 = 3'h0;
  wire [0:0] v_3883_0;
  wire [0:0] v_3884_0;
  wire [0:0] v_3885_0;
  wire [2:0] v_3886_0;
  wire [2:0] v_3887_0;
  wire [2:0] v_3888_0;
  reg [2:0] v_3889_0 = 3'h0;
  wire [0:0] v_3890_0;
  wire [0:0] v_3891_0;
  wire [0:0] v_3892_0;
  wire [2:0] v_3893_0;
  wire [2:0] v_3894_0;
  wire [2:0] v_3895_0;
  reg [2:0] v_3896_0 = 3'h0;
  wire [0:0] v_3897_0;
  wire [0:0] v_3898_0;
  wire [0:0] v_3899_0;
  wire [2:0] v_3900_0;
  wire [2:0] v_3901_0;
  wire [2:0] v_3902_0;
  reg [2:0] v_3903_0 = 3'h0;
  wire [0:0] v_3904_0;
  wire [0:0] v_3905_0;
  wire [0:0] v_3906_0;
  wire [2:0] v_3907_0;
  wire [2:0] v_3908_0;
  wire [2:0] v_3909_0;
  reg [2:0] v_3910_0 = 3'h0;
  wire [0:0] v_3911_0;
  wire [0:0] v_3912_0;
  wire [0:0] v_3913_0;
  wire [2:0] v_3914_0;
  wire [2:0] v_3915_0;
  wire [2:0] v_3916_0;
  reg [2:0] v_3917_0 = 3'h0;
  wire [0:0] v_3918_0;
  wire [0:0] v_3919_0;
  wire [0:0] v_3920_0;
  wire [2:0] v_3921_0;
  wire [2:0] v_3922_0;
  wire [2:0] v_3923_0;
  reg [2:0] v_3924_0 = 3'h0;
  wire [0:0] v_3925_0;
  wire [0:0] v_3926_0;
  wire [0:0] v_3927_0;
  wire [2:0] v_3928_0;
  wire [2:0] v_3929_0;
  wire [2:0] v_3930_0;
  reg [2:0] v_3931_0 = 3'h0;
  wire [0:0] v_3932_0;
  wire [0:0] v_3933_0;
  wire [0:0] v_3934_0;
  wire [2:0] v_3935_0;
  wire [2:0] v_3936_0;
  wire [2:0] v_3937_0;
  reg [2:0] v_3938_0 = 3'h0;
  wire [0:0] v_3939_0;
  wire [0:0] v_3940_0;
  wire [0:0] v_3941_0;
  wire [2:0] v_3942_0;
  wire [2:0] v_3943_0;
  wire [2:0] v_3944_0;
  reg [2:0] v_3945_0 = 3'h0;
  wire [0:0] v_3946_0;
  wire [0:0] v_3947_0;
  wire [0:0] v_3948_0;
  wire [2:0] v_3949_0;
  wire [2:0] v_3950_0;
  wire [2:0] v_3951_0;
  reg [2:0] v_3952_0 = 3'h0;
  wire [0:0] v_3953_0;
  wire [0:0] v_3954_0;
  wire [0:0] v_3955_0;
  wire [2:0] v_3956_0;
  wire [2:0] v_3957_0;
  wire [2:0] v_3958_0;
  reg [2:0] v_3959_0 = 3'h0;
  wire [0:0] v_3960_0;
  wire [0:0] v_3961_0;
  wire [0:0] v_3962_0;
  wire [2:0] v_3963_0;
  wire [2:0] v_3964_0;
  wire [2:0] v_3965_0;
  reg [2:0] v_3966_0 = 3'h0;
  wire [0:0] v_3967_0;
  wire [0:0] v_3968_0;
  wire [0:0] v_3969_0;
  wire [2:0] v_3970_0;
  wire [2:0] v_3971_0;
  wire [2:0] v_3972_0;
  reg [2:0] v_3973_0 = 3'h0;
  wire [0:0] v_3974_0;
  wire [0:0] v_3975_0;
  wire [0:0] v_3976_0;
  wire [2:0] v_3977_0;
  wire [2:0] v_3978_0;
  wire [2:0] v_3979_0;
  reg [2:0] v_3980_0 = 3'h0;
  wire [0:0] v_3981_0;
  wire [0:0] v_3982_0;
  wire [0:0] v_3983_0;
  wire [2:0] v_3984_0;
  wire [2:0] v_3985_0;
  wire [2:0] v_3986_0;
  reg [2:0] v_3987_0 = 3'h0;
  wire [0:0] v_3988_0;
  wire [0:0] v_3989_0;
  wire [0:0] v_3990_0;
  wire [2:0] v_3991_0;
  wire [2:0] v_3992_0;
  wire [2:0] v_3993_0;
  reg [2:0] v_3994_0 = 3'h0;
  wire [0:0] v_3995_0;
  wire [0:0] v_3996_0;
  wire [0:0] v_3997_0;
  wire [2:0] v_3998_0;
  wire [2:0] v_3999_0;
  wire [2:0] v_4000_0;
  reg [2:0] v_4001_0 = 3'h0;
  wire [0:0] v_4002_0;
  wire [0:0] v_4003_0;
  wire [0:0] v_4004_0;
  wire [2:0] v_4005_0;
  wire [2:0] v_4006_0;
  wire [2:0] v_4007_0;
  reg [2:0] v_4008_0 = 3'h0;
  wire [0:0] v_4009_0;
  wire [0:0] v_4010_0;
  wire [0:0] v_4011_0;
  wire [2:0] v_4012_0;
  wire [2:0] v_4013_0;
  wire [2:0] v_4014_0;
  reg [2:0] v_4015_0 = 3'h0;
  wire [0:0] v_4016_0;
  wire [0:0] v_4017_0;
  wire [0:0] v_4018_0;
  wire [2:0] v_4019_0;
  wire [2:0] v_4020_0;
  wire [2:0] v_4021_0;
  reg [2:0] v_4022_0 = 3'h0;
  wire [0:0] v_4023_0;
  wire [0:0] v_4024_0;
  wire [0:0] v_4025_0;
  wire [2:0] v_4026_0;
  wire [2:0] v_4027_0;
  wire [2:0] v_4028_0;
  reg [2:0] v_4029_0 = 3'h0;
  wire [0:0] v_4030_0;
  wire [0:0] v_4031_0;
  wire [0:0] v_4032_0;
  wire [2:0] v_4033_0;
  wire [2:0] v_4034_0;
  wire [2:0] v_4035_0;
  reg [2:0] v_4036_0 = 3'h0;
  wire [0:0] v_4037_0;
  wire [0:0] v_4038_0;
  wire [0:0] v_4039_0;
  wire [2:0] v_4040_0;
  wire [2:0] v_4041_0;
  wire [2:0] v_4042_0;
  reg [2:0] v_4043_0 = 3'h0;
  wire [0:0] v_4044_0;
  wire [0:0] v_4045_0;
  wire [0:0] v_4046_0;
  wire [2:0] v_4047_0;
  wire [2:0] v_4048_0;
  wire [2:0] v_4049_0;
  reg [2:0] v_4050_0 = 3'h0;
  wire [0:0] v_4051_0;
  wire [0:0] v_4052_0;
  wire [0:0] v_4053_0;
  wire [2:0] v_4054_0;
  wire [2:0] v_4055_0;
  wire [2:0] v_4056_0;
  reg [2:0] v_4057_0 = 3'h0;
  wire [0:0] v_4058_0;
  wire [0:0] v_4059_0;
  wire [0:0] v_4060_0;
  wire [2:0] v_4061_0;
  wire [2:0] v_4062_0;
  wire [2:0] v_4063_0;
  reg [2:0] v_4064_0 = 3'h0;
  wire [0:0] v_4065_0;
  wire [0:0] v_4066_0;
  wire [0:0] v_4067_0;
  wire [2:0] v_4068_0;
  wire [2:0] v_4069_0;
  wire [2:0] v_4070_0;
  reg [2:0] v_4071_0 = 3'h0;
  wire [0:0] v_4072_0;
  wire [0:0] v_4073_0;
  wire [0:0] v_4074_0;
  wire [2:0] v_4075_0;
  wire [2:0] v_4076_0;
  wire [2:0] v_4077_0;
  reg [2:0] v_4078_0 = 3'h0;
  wire [0:0] v_4079_0;
  wire [0:0] v_4080_0;
  wire [0:0] v_4081_0;
  wire [2:0] v_4082_0;
  wire [2:0] v_4083_0;
  wire [2:0] v_4084_0;
  reg [2:0] v_4085_0 = 3'h0;
  wire [0:0] v_4086_0;
  wire [0:0] v_4087_0;
  wire [0:0] v_4088_0;
  wire [2:0] v_4089_0;
  wire [2:0] v_4090_0;
  wire [2:0] v_4091_0;
  reg [2:0] v_4092_0 = 3'h0;
  wire [0:0] v_4093_0;
  wire [0:0] v_4094_0;
  wire [0:0] v_4095_0;
  wire [2:0] v_4096_0;
  wire [2:0] v_4097_0;
  wire [2:0] v_4098_0;
  reg [2:0] v_4099_0 = 3'h0;
  wire [0:0] v_4100_0;
  wire [0:0] v_4101_0;
  wire [0:0] v_4102_0;
  wire [2:0] v_4103_0;
  wire [2:0] v_4104_0;
  wire [2:0] v_4105_0;
  reg [2:0] v_4106_0 = 3'h0;
  wire [0:0] v_4107_0;
  wire [0:0] v_4108_0;
  wire [0:0] v_4109_0;
  wire [2:0] v_4110_0;
  wire [2:0] v_4111_0;
  wire [2:0] v_4112_0;
  reg [2:0] v_4113_0 = 3'h0;
  wire [0:0] v_4114_0;
  wire [0:0] v_4115_0;
  wire [0:0] v_4116_0;
  wire [2:0] v_4117_0;
  wire [2:0] v_4118_0;
  wire [2:0] v_4119_0;
  reg [2:0] v_4120_0 = 3'h0;
  wire [0:0] v_4121_0;
  wire [0:0] v_4122_0;
  wire [0:0] v_4123_0;
  wire [2:0] v_4124_0;
  wire [2:0] v_4125_0;
  wire [2:0] v_4126_0;
  reg [2:0] v_4127_0 = 3'h0;
  wire [0:0] v_4128_0;
  wire [0:0] v_4129_0;
  wire [0:0] v_4130_0;
  wire [2:0] v_4131_0;
  wire [2:0] v_4132_0;
  wire [2:0] v_4133_0;
  reg [2:0] v_4134_0 = 3'h0;
  wire [0:0] v_4135_0;
  wire [0:0] v_4136_0;
  wire [0:0] v_4137_0;
  wire [2:0] v_4138_0;
  wire [2:0] v_4139_0;
  wire [2:0] v_4140_0;
  reg [2:0] v_4141_0 = 3'h0;
  wire [0:0] v_4142_0;
  wire [0:0] v_4143_0;
  wire [0:0] v_4144_0;
  wire [2:0] v_4145_0;
  wire [2:0] v_4146_0;
  wire [2:0] v_4147_0;
  reg [2:0] v_4148_0 = 3'h0;
  wire [0:0] v_4149_0;
  wire [0:0] v_4150_0;
  wire [0:0] v_4151_0;
  wire [2:0] v_4152_0;
  wire [2:0] v_4153_0;
  wire [2:0] v_4154_0;
  reg [2:0] v_4155_0 = 3'h0;
  wire [0:0] v_4156_0;
  wire [0:0] v_4157_0;
  wire [0:0] v_4158_0;
  wire [2:0] v_4159_0;
  wire [2:0] v_4160_0;
  wire [2:0] v_4161_0;
  reg [2:0] v_4162_0 = 3'h0;
  wire [0:0] v_4163_0;
  wire [0:0] v_4164_0;
  wire [0:0] v_4165_0;
  wire [2:0] v_4166_0;
  wire [2:0] v_4167_0;
  wire [2:0] v_4168_0;
  reg [2:0] v_4169_0 = 3'h0;
  wire [0:0] v_4170_0;
  wire [0:0] v_4171_0;
  wire [0:0] v_4172_0;
  wire [2:0] v_4173_0;
  wire [2:0] v_4174_0;
  wire [2:0] v_4175_0;
  reg [2:0] v_4176_0 = 3'h0;
  wire [0:0] v_4177_0;
  wire [0:0] v_4178_0;
  wire [0:0] v_4179_0;
  wire [2:0] v_4180_0;
  wire [2:0] v_4181_0;
  wire [2:0] v_4182_0;
  reg [2:0] v_4183_0 = 3'h0;
  wire [0:0] v_4184_0;
  wire [0:0] v_4185_0;
  wire [0:0] v_4186_0;
  wire [2:0] v_4187_0;
  wire [2:0] v_4188_0;
  wire [2:0] v_4189_0;
  reg [2:0] v_4190_0 = 3'h0;
  wire [0:0] v_4191_0;
  wire [0:0] v_4192_0;
  wire [0:0] v_4193_0;
  wire [2:0] v_4194_0;
  wire [2:0] v_4195_0;
  wire [2:0] v_4196_0;
  reg [2:0] v_4197_0 = 3'h0;
  wire [0:0] v_4198_0;
  wire [0:0] v_4199_0;
  wire [0:0] v_4200_0;
  wire [2:0] v_4201_0;
  wire [2:0] v_4202_0;
  wire [2:0] v_4203_0;
  reg [2:0] v_4204_0 = 3'h0;
  wire [0:0] v_4205_0;
  wire [0:0] v_4206_0;
  wire [0:0] v_4207_0;
  wire [2:0] v_4208_0;
  wire [2:0] v_4209_0;
  wire [2:0] v_4210_0;
  reg [2:0] v_4211_0 = 3'h0;
  wire [0:0] v_4212_0;
  wire [0:0] v_4213_0;
  wire [0:0] v_4214_0;
  wire [2:0] v_4215_0;
  wire [2:0] v_4216_0;
  wire [2:0] v_4217_0;
  reg [2:0] v_4218_0 = 3'h0;
  wire [0:0] v_4219_0;
  wire [0:0] v_4220_0;
  wire [0:0] v_4221_0;
  wire [2:0] v_4222_0;
  wire [2:0] v_4223_0;
  wire [2:0] v_4224_0;
  reg [2:0] v_4225_0 = 3'h0;
  wire [0:0] v_4226_0;
  wire [0:0] v_4227_0;
  wire [0:0] v_4228_0;
  wire [2:0] v_4229_0;
  wire [2:0] v_4230_0;
  wire [2:0] v_4231_0;
  reg [2:0] v_4232_0 = 3'h0;
  wire [0:0] v_4233_0;
  wire [0:0] v_4234_0;
  wire [0:0] v_4235_0;
  wire [2:0] v_4236_0;
  wire [2:0] v_4237_0;
  wire [2:0] v_4238_0;
  reg [2:0] v_4239_0 = 3'h0;
  wire [0:0] v_4240_0;
  wire [0:0] v_4241_0;
  wire [0:0] v_4242_0;
  wire [2:0] v_4243_0;
  wire [2:0] v_4244_0;
  wire [2:0] v_4245_0;
  reg [2:0] v_4246_0 = 3'h0;
  wire [0:0] v_4247_0;
  wire [0:0] v_4248_0;
  wire [0:0] v_4249_0;
  wire [2:0] v_4250_0;
  wire [2:0] v_4251_0;
  wire [2:0] v_4252_0;
  reg [2:0] v_4253_0 = 3'h0;
  wire [0:0] v_4254_0;
  wire [0:0] v_4255_0;
  wire [0:0] v_4256_0;
  wire [2:0] v_4257_0;
  wire [2:0] v_4258_0;
  wire [2:0] v_4259_0;
  reg [2:0] v_4260_0 = 3'h0;
  wire [0:0] v_4261_0;
  wire [0:0] v_4262_0;
  wire [0:0] v_4263_0;
  wire [2:0] v_4264_0;
  wire [2:0] v_4265_0;
  wire [2:0] v_4266_0;
  reg [2:0] v_4267_0 = 3'h0;
  wire [0:0] v_4268_0;
  wire [0:0] v_4269_0;
  wire [0:0] v_4270_0;
  wire [2:0] v_4271_0;
  wire [2:0] v_4272_0;
  wire [2:0] v_4273_0;
  reg [2:0] v_4274_0 = 3'h0;
  wire [0:0] v_4275_0;
  wire [0:0] v_4276_0;
  wire [0:0] v_4277_0;
  wire [2:0] v_4278_0;
  wire [2:0] v_4279_0;
  wire [2:0] v_4280_0;
  reg [2:0] v_4281_0 = 3'h0;
  wire [0:0] v_4282_0;
  wire [0:0] v_4283_0;
  wire [0:0] v_4284_0;
  wire [2:0] v_4285_0;
  wire [2:0] v_4286_0;
  wire [2:0] v_4287_0;
  reg [2:0] v_4288_0 = 3'h0;
  wire [0:0] v_4289_0;
  wire [0:0] v_4290_0;
  wire [0:0] v_4291_0;
  wire [2:0] v_4292_0;
  wire [2:0] v_4293_0;
  wire [2:0] v_4294_0;
  reg [2:0] v_4295_0 = 3'h0;
  wire [0:0] v_4296_0;
  wire [0:0] v_4297_0;
  wire [0:0] v_4298_0;
  wire [2:0] v_4299_0;
  wire [2:0] v_4300_0;
  wire [2:0] v_4301_0;
  reg [2:0] v_4302_0 = 3'h0;
  wire [0:0] v_4303_0;
  wire [0:0] v_4304_0;
  wire [0:0] v_4305_0;
  wire [2:0] v_4306_0;
  wire [2:0] v_4307_0;
  wire [2:0] v_4308_0;
  reg [2:0] v_4309_0 = 3'h0;
  wire [0:0] v_4310_0;
  wire [0:0] v_4311_0;
  wire [0:0] v_4312_0;
  wire [2:0] v_4313_0;
  wire [2:0] v_4314_0;
  wire [2:0] v_4315_0;
  reg [2:0] v_4316_0 = 3'h0;
  wire [0:0] v_4317_0;
  wire [0:0] v_4318_0;
  wire [0:0] v_4319_0;
  wire [2:0] v_4320_0;
  wire [2:0] v_4321_0;
  wire [2:0] v_4322_0;
  reg [2:0] v_4323_0 = 3'h0;
  wire [0:0] v_4324_0;
  wire [0:0] v_4325_0;
  wire [0:0] v_4326_0;
  wire [2:0] v_4327_0;
  wire [2:0] v_4328_0;
  wire [2:0] v_4329_0;
  reg [2:0] v_4330_0 = 3'h0;
  wire [0:0] v_4331_0;
  wire [0:0] v_4332_0;
  wire [0:0] v_4333_0;
  wire [2:0] v_4334_0;
  wire [2:0] v_4335_0;
  wire [2:0] v_4336_0;
  reg [2:0] v_4337_0 = 3'h0;
  wire [0:0] v_4338_0;
  wire [0:0] v_4339_0;
  wire [0:0] v_4340_0;
  wire [2:0] v_4341_0;
  wire [2:0] v_4342_0;
  wire [2:0] v_4343_0;
  reg [2:0] v_4344_0 = 3'h0;
  wire [0:0] v_4345_0;
  wire [0:0] v_4346_0;
  wire [0:0] v_4347_0;
  wire [2:0] v_4348_0;
  wire [2:0] v_4349_0;
  wire [2:0] v_4350_0;
  reg [2:0] v_4351_0 = 3'h0;
  wire [0:0] v_4352_0;
  wire [0:0] v_4353_0;
  wire [0:0] v_4354_0;
  wire [2:0] v_4355_0;
  wire [2:0] v_4356_0;
  wire [2:0] v_4357_0;
  reg [2:0] v_4358_0 = 3'h0;
  wire [0:0] v_4359_0;
  wire [0:0] v_4360_0;
  wire [0:0] v_4361_0;
  wire [2:0] v_4362_0;
  wire [2:0] v_4363_0;
  wire [2:0] v_4364_0;
  reg [2:0] v_4365_0 = 3'h0;
  wire [0:0] v_4366_0;
  wire [0:0] v_4367_0;
  wire [0:0] v_4368_0;
  wire [2:0] v_4369_0;
  wire [2:0] v_4370_0;
  wire [2:0] v_4371_0;
  reg [2:0] v_4372_0 = 3'h0;
  wire [0:0] v_4373_0;
  wire [0:0] v_4374_0;
  wire [0:0] v_4375_0;
  wire [2:0] v_4376_0;
  wire [2:0] v_4377_0;
  wire [2:0] v_4378_0;
  reg [2:0] v_4379_0 = 3'h0;
  wire [0:0] v_4380_0;
  wire [0:0] v_4381_0;
  wire [0:0] v_4382_0;
  wire [2:0] v_4383_0;
  wire [2:0] v_4384_0;
  wire [2:0] v_4385_0;
  reg [2:0] v_4386_0 = 3'h0;
  wire [0:0] v_4387_0;
  wire [0:0] v_4388_0;
  wire [0:0] v_4389_0;
  wire [2:0] v_4390_0;
  wire [2:0] v_4391_0;
  wire [2:0] v_4392_0;
  reg [2:0] v_4393_0 = 3'h0;
  wire [0:0] v_4394_0;
  wire [0:0] v_4395_0;
  wire [0:0] v_4396_0;
  wire [2:0] v_4397_0;
  wire [2:0] v_4398_0;
  wire [2:0] v_4399_0;
  reg [2:0] v_4400_0 = 3'h0;
  wire [0:0] v_4401_0;
  wire [0:0] v_4402_0;
  wire [0:0] v_4403_0;
  wire [2:0] v_4404_0;
  wire [2:0] v_4405_0;
  wire [2:0] v_4406_0;
  reg [2:0] v_4407_0 = 3'h0;
  wire [0:0] v_4408_0;
  wire [0:0] v_4409_0;
  wire [0:0] v_4410_0;
  wire [2:0] v_4411_0;
  wire [2:0] v_4412_0;
  wire [2:0] v_4413_0;
  reg [2:0] v_4414_0 = 3'h0;
  wire [0:0] v_4415_0;
  wire [0:0] v_4416_0;
  wire [0:0] v_4417_0;
  wire [2:0] v_4418_0;
  wire [2:0] v_4419_0;
  wire [2:0] v_4420_0;
  reg [2:0] v_4421_0 = 3'h0;
  wire [0:0] v_4422_0;
  wire [0:0] v_4423_0;
  wire [0:0] v_4424_0;
  wire [2:0] v_4425_0;
  wire [2:0] v_4426_0;
  wire [2:0] v_4427_0;
  reg [2:0] v_4428_0 = 3'h0;
  wire [0:0] v_4429_0;
  wire [0:0] v_4430_0;
  wire [0:0] v_4431_0;
  wire [2:0] v_4432_0;
  wire [2:0] v_4433_0;
  wire [2:0] v_4434_0;
  reg [2:0] v_4435_0 = 3'h0;
  wire [0:0] v_4436_0;
  wire [0:0] v_4437_0;
  wire [0:0] v_4438_0;
  wire [2:0] v_4439_0;
  wire [2:0] v_4440_0;
  wire [2:0] v_4441_0;
  reg [2:0] v_4442_0 = 3'h0;
  wire [0:0] v_4443_0;
  wire [0:0] v_4444_0;
  wire [0:0] v_4445_0;
  wire [2:0] v_4446_0;
  wire [2:0] v_4447_0;
  wire [2:0] v_4448_0;
  reg [2:0] v_4449_0 = 3'h0;
  wire [0:0] v_4450_0;
  wire [0:0] v_4451_0;
  wire [0:0] v_4452_0;
  wire [2:0] v_4453_0;
  wire [2:0] v_4454_0;
  wire [2:0] v_4455_0;
  reg [2:0] v_4456_0 = 3'h0;
  wire [0:0] v_4457_0;
  wire [0:0] v_4458_0;
  wire [0:0] v_4459_0;
  wire [2:0] v_4460_0;
  wire [2:0] v_4461_0;
  wire [2:0] v_4462_0;
  reg [2:0] v_4463_0 = 3'h0;
  wire [0:0] v_4464_0;
  wire [0:0] v_4465_0;
  wire [0:0] v_4466_0;
  wire [2:0] v_4467_0;
  wire [2:0] v_4468_0;
  wire [2:0] v_4469_0;
  reg [2:0] v_4470_0 = 3'h0;
  wire [0:0] v_4471_0;
  wire [0:0] v_4472_0;
  wire [0:0] v_4473_0;
  wire [2:0] v_4474_0;
  wire [2:0] v_4475_0;
  wire [2:0] v_4476_0;
  reg [2:0] v_4477_0 = 3'h0;
  wire [0:0] v_4478_0;
  wire [0:0] v_4479_0;
  wire [0:0] v_4480_0;
  wire [2:0] v_4481_0;
  wire [2:0] v_4482_0;
  wire [2:0] v_4483_0;
  reg [2:0] v_4484_0 = 3'h0;
  wire [0:0] v_4485_0;
  wire [0:0] v_4486_0;
  wire [0:0] v_4487_0;
  wire [2:0] v_4488_0;
  wire [2:0] v_4489_0;
  wire [2:0] v_4490_0;
  reg [2:0] v_4491_0 = 3'h0;
  wire [0:0] v_4492_0;
  wire [0:0] v_4493_0;
  wire [0:0] v_4494_0;
  wire [2:0] v_4495_0;
  wire [2:0] v_4496_0;
  wire [2:0] v_4497_0;
  reg [2:0] v_4498_0 = 3'h0;
  wire [0:0] v_4499_0;
  wire [0:0] v_4500_0;
  wire [0:0] v_4501_0;
  wire [2:0] v_4502_0;
  wire [2:0] v_4503_0;
  wire [2:0] v_4504_0;
  reg [2:0] v_4505_0 = 3'h0;
  wire [0:0] v_4506_0;
  wire [0:0] v_4507_0;
  wire [0:0] v_4508_0;
  wire [2:0] v_4509_0;
  wire [2:0] v_4510_0;
  wire [2:0] v_4511_0;
  reg [2:0] v_4512_0 = 3'h0;
  wire [0:0] v_4513_0;
  wire [0:0] v_4514_0;
  wire [0:0] v_4515_0;
  wire [2:0] v_4516_0;
  wire [2:0] v_4517_0;
  wire [2:0] v_4518_0;
  reg [2:0] v_4519_0 = 3'h0;
  wire [0:0] v_4520_0;
  wire [0:0] v_4521_0;
  wire [0:0] v_4522_0;
  wire [2:0] v_4523_0;
  wire [2:0] v_4524_0;
  wire [2:0] v_4525_0;
  reg [2:0] v_4526_0 = 3'h0;
  wire [0:0] v_4527_0;
  wire [0:0] v_4528_0;
  wire [0:0] v_4529_0;
  wire [2:0] v_4530_0;
  wire [2:0] v_4531_0;
  wire [2:0] v_4532_0;
  reg [2:0] v_4533_0 = 3'h0;
  wire [0:0] v_4534_0;
  wire [0:0] v_4535_0;
  wire [0:0] v_4536_0;
  wire [2:0] v_4537_0;
  wire [2:0] v_4538_0;
  wire [2:0] v_4539_0;
  reg [2:0] v_4540_0 = 3'h0;
  wire [0:0] v_4541_0;
  wire [0:0] v_4542_0;
  wire [0:0] v_4543_0;
  wire [2:0] v_4544_0;
  wire [2:0] v_4545_0;
  wire [2:0] v_4546_0;
  reg [2:0] v_4547_0 = 3'h0;
  wire [0:0] v_4548_0;
  wire [0:0] v_4549_0;
  wire [0:0] v_4550_0;
  wire [2:0] v_4551_0;
  wire [2:0] v_4552_0;
  wire [2:0] v_4553_0;
  reg [2:0] v_4554_0 = 3'h0;
  wire [0:0] v_4555_0;
  wire [0:0] v_4556_0;
  wire [0:0] v_4557_0;
  wire [2:0] v_4558_0;
  wire [2:0] v_4559_0;
  wire [2:0] v_4560_0;
  reg [2:0] v_4561_0 = 3'h0;
  wire [0:0] v_4562_0;
  wire [0:0] v_4563_0;
  wire [0:0] v_4564_0;
  wire [2:0] v_4565_0;
  wire [2:0] v_4566_0;
  wire [2:0] v_4567_0;
  reg [2:0] v_4568_0 = 3'h0;
  wire [0:0] v_4569_0;
  wire [0:0] v_4570_0;
  wire [0:0] v_4571_0;
  wire [2:0] v_4572_0;
  wire [2:0] v_4573_0;
  wire [2:0] v_4574_0;
  reg [2:0] v_4575_0 = 3'h0;
  wire [0:0] v_4576_0;
  wire [0:0] v_4577_0;
  wire [0:0] v_4578_0;
  wire [2:0] v_4579_0;
  wire [2:0] v_4580_0;
  wire [2:0] v_4581_0;
  reg [2:0] v_4582_0 = 3'h0;
  wire [0:0] v_4583_0;
  wire [0:0] v_4584_0;
  wire [0:0] v_4585_0;
  wire [2:0] v_4586_0;
  wire [2:0] v_4587_0;
  wire [2:0] v_4588_0;
  reg [2:0] v_4589_0 = 3'h0;
  wire [0:0] v_4590_0;
  wire [0:0] v_4591_0;
  wire [0:0] v_4592_0;
  wire [2:0] v_4593_0;
  wire [2:0] v_4594_0;
  wire [2:0] v_4595_0;
  reg [2:0] v_4596_0 = 3'h0;
  wire [0:0] v_4597_0;
  wire [0:0] v_4598_0;
  wire [0:0] v_4599_0;
  wire [2:0] v_4600_0;
  wire [2:0] v_4601_0;
  wire [2:0] v_4602_0;
  reg [2:0] v_4603_0 = 3'h0;
  wire [0:0] v_4604_0;
  wire [0:0] v_4605_0;
  wire [0:0] v_4606_0;
  wire [2:0] v_4607_0;
  wire [2:0] v_4608_0;
  wire [2:0] v_4609_0;
  reg [2:0] v_4610_0 = 3'h0;
  wire [0:0] v_4611_0;
  wire [0:0] v_4612_0;
  wire [0:0] v_4613_0;
  wire [2:0] v_4614_0;
  wire [2:0] v_4615_0;
  wire [2:0] v_4616_0;
  reg [2:0] v_4617_0 = 3'h0;
  wire [0:0] v_4618_0;
  wire [0:0] v_4619_0;
  wire [0:0] v_4620_0;
  wire [2:0] v_4621_0;
  wire [2:0] v_4622_0;
  wire [2:0] v_4623_0;
  reg [2:0] v_4624_0 = 3'h0;
  wire [0:0] v_4625_0;
  wire [0:0] v_4626_0;
  wire [0:0] v_4627_0;
  wire [2:0] v_4628_0;
  wire [2:0] v_4629_0;
  wire [2:0] v_4630_0;
  reg [2:0] v_4631_0 = 3'h0;
  wire [0:0] v_4632_0;
  wire [0:0] v_4633_0;
  wire [0:0] v_4634_0;
  wire [2:0] v_4635_0;
  wire [2:0] v_4636_0;
  wire [2:0] v_4637_0;
  reg [2:0] v_4638_0 = 3'h0;
  wire [0:0] v_4639_0;
  wire [0:0] v_4640_0;
  wire [0:0] v_4641_0;
  wire [2:0] v_4642_0;
  wire [2:0] v_4643_0;
  wire [2:0] v_4644_0;
  reg [2:0] v_4645_0 = 3'h0;
  wire [0:0] v_4646_0;
  wire [0:0] v_4647_0;
  wire [0:0] v_4648_0;
  wire [2:0] v_4649_0;
  wire [2:0] v_4650_0;
  wire [2:0] v_4651_0;
  reg [2:0] v_4652_0 = 3'h0;
  wire [0:0] v_4653_0;
  wire [0:0] v_4654_0;
  wire [0:0] v_4655_0;
  wire [2:0] v_4656_0;
  wire [2:0] v_4657_0;
  wire [2:0] v_4658_0;
  reg [2:0] v_4659_0 = 3'h0;
  wire [0:0] v_4660_0;
  wire [0:0] v_4661_0;
  wire [0:0] v_4662_0;
  wire [2:0] v_4663_0;
  wire [2:0] v_4664_0;
  wire [2:0] v_4665_0;
  reg [2:0] v_4666_0 = 3'h0;
  wire [0:0] v_4667_0;
  wire [0:0] v_4668_0;
  wire [0:0] v_4669_0;
  wire [2:0] v_4670_0;
  wire [2:0] v_4671_0;
  wire [2:0] v_4672_0;
  reg [2:0] v_4673_0 = 3'h0;
  wire [0:0] v_4674_0;
  wire [0:0] v_4675_0;
  wire [0:0] v_4676_0;
  wire [2:0] v_4677_0;
  wire [2:0] v_4678_0;
  wire [2:0] v_4679_0;
  reg [2:0] v_4680_0 = 3'h0;
  wire [0:0] v_4681_0;
  wire [0:0] v_4682_0;
  wire [0:0] v_4683_0;
  wire [2:0] v_4684_0;
  wire [2:0] v_4685_0;
  wire [2:0] v_4686_0;
  reg [2:0] v_4687_0 = 3'h0;
  wire [0:0] v_4688_0;
  wire [0:0] v_4689_0;
  wire [0:0] v_4690_0;
  wire [2:0] v_4691_0;
  wire [2:0] v_4692_0;
  wire [2:0] v_4693_0;
  reg [2:0] v_4694_0 = 3'h0;
  wire [0:0] v_4695_0;
  wire [0:0] v_4696_0;
  wire [0:0] v_4697_0;
  wire [2:0] v_4698_0;
  wire [2:0] v_4699_0;
  wire [2:0] v_4700_0;
  reg [2:0] v_4701_0 = 3'h0;
  wire [0:0] v_4702_0;
  wire [0:0] v_4703_0;
  wire [0:0] v_4704_0;
  wire [2:0] v_4705_0;
  wire [2:0] v_4706_0;
  wire [2:0] v_4707_0;
  reg [2:0] v_4708_0 = 3'h0;
  wire [0:0] v_4709_0;
  wire [0:0] v_4710_0;
  wire [0:0] v_4711_0;
  wire [2:0] v_4712_0;
  wire [2:0] v_4713_0;
  wire [2:0] v_4714_0;
  reg [2:0] v_4715_0 = 3'h0;
  wire [0:0] v_4716_0;
  wire [0:0] v_4717_0;
  wire [0:0] v_4718_0;
  wire [2:0] v_4719_0;
  wire [2:0] v_4720_0;
  wire [2:0] v_4721_0;
  reg [2:0] v_4722_0 = 3'h0;
  wire [0:0] v_4723_0;
  wire [0:0] v_4724_0;
  wire [0:0] v_4725_0;
  wire [2:0] v_4726_0;
  wire [2:0] v_4727_0;
  wire [2:0] v_4728_0;
  reg [2:0] v_4729_0 = 3'h0;
  wire [0:0] v_4730_0;
  wire [0:0] v_4731_0;
  wire [0:0] v_4732_0;
  wire [2:0] v_4733_0;
  wire [2:0] v_4734_0;
  wire [2:0] v_4735_0;
  reg [2:0] v_4736_0 = 3'h0;
  wire [0:0] v_4737_0;
  wire [0:0] v_4738_0;
  wire [0:0] v_4739_0;
  wire [2:0] v_4740_0;
  wire [2:0] v_4741_0;
  wire [2:0] v_4742_0;
  reg [2:0] v_4743_0 = 3'h0;
  wire [0:0] v_4744_0;
  wire [0:0] v_4745_0;
  wire [0:0] v_4746_0;
  wire [2:0] v_4747_0;
  wire [2:0] v_4748_0;
  wire [2:0] v_4749_0;
  reg [2:0] v_4750_0 = 3'h0;
  wire [0:0] v_4751_0;
  wire [0:0] v_4752_0;
  wire [0:0] v_4753_0;
  wire [2:0] v_4754_0;
  wire [2:0] v_4755_0;
  wire [2:0] v_4756_0;
  reg [2:0] v_4757_0 = 3'h0;
  wire [0:0] v_4758_0;
  wire [0:0] v_4759_0;
  wire [0:0] v_4760_0;
  wire [2:0] v_4761_0;
  wire [2:0] v_4762_0;
  wire [2:0] v_4763_0;
  reg [2:0] v_4764_0 = 3'h0;
  wire [0:0] v_4765_0;
  wire [0:0] v_4766_0;
  wire [0:0] v_4767_0;
  wire [2:0] v_4768_0;
  wire [2:0] v_4769_0;
  wire [2:0] v_4770_0;
  reg [2:0] v_4771_0 = 3'h0;
  wire [0:0] v_4772_0;
  wire [0:0] v_4773_0;
  wire [0:0] v_4774_0;
  wire [2:0] v_4775_0;
  wire [2:0] v_4776_0;
  wire [2:0] v_4777_0;
  reg [2:0] v_4778_0 = 3'h0;
  wire [0:0] v_4779_0;
  wire [0:0] v_4780_0;
  wire [0:0] v_4781_0;
  wire [2:0] v_4782_0;
  wire [2:0] v_4783_0;
  wire [2:0] v_4784_0;
  reg [2:0] v_4785_0 = 3'h0;
  wire [0:0] v_4786_0;
  wire [0:0] v_4787_0;
  wire [0:0] v_4788_0;
  wire [2:0] v_4789_0;
  wire [2:0] v_4790_0;
  wire [2:0] v_4791_0;
  reg [2:0] v_4792_0 = 3'h0;
  wire [0:0] v_4793_0;
  wire [0:0] v_4794_0;
  wire [0:0] v_4795_0;
  wire [2:0] v_4796_0;
  wire [2:0] v_4797_0;
  wire [2:0] v_4798_0;
  reg [2:0] v_4799_0 = 3'h0;
  wire [0:0] v_4800_0;
  wire [0:0] v_4801_0;
  wire [0:0] v_4802_0;
  wire [2:0] v_4803_0;
  wire [2:0] v_4804_0;
  wire [2:0] v_4805_0;
  reg [2:0] v_4806_0 = 3'h0;
  wire [0:0] v_4807_0;
  wire [0:0] v_4808_0;
  wire [0:0] v_4809_0;
  wire [2:0] v_4810_0;
  wire [2:0] v_4811_0;
  wire [2:0] v_4812_0;
  reg [2:0] v_4813_0 = 3'h0;
  wire [0:0] v_4814_0;
  wire [0:0] v_4815_0;
  wire [0:0] v_4816_0;
  wire [2:0] v_4817_0;
  wire [2:0] v_4818_0;
  wire [2:0] v_4819_0;
  reg [2:0] v_4820_0 = 3'h0;
  wire [0:0] v_4821_0;
  wire [0:0] v_4822_0;
  wire [0:0] v_4823_0;
  wire [2:0] v_4824_0;
  wire [2:0] v_4825_0;
  wire [2:0] v_4826_0;
  reg [2:0] v_4827_0 = 3'h0;
  wire [0:0] v_4828_0;
  wire [0:0] v_4829_0;
  wire [0:0] v_4830_0;
  wire [2:0] v_4831_0;
  wire [2:0] v_4832_0;
  wire [2:0] v_4833_0;
  reg [2:0] v_4834_0 = 3'h0;
  wire [0:0] v_4835_0;
  wire [0:0] v_4836_0;
  wire [0:0] v_4837_0;
  wire [2:0] v_4838_0;
  wire [2:0] v_4839_0;
  wire [2:0] v_4840_0;
  reg [2:0] v_4841_0 = 3'h0;
  wire [0:0] v_4842_0;
  wire [0:0] v_4843_0;
  wire [0:0] v_4844_0;
  wire [2:0] v_4845_0;
  wire [2:0] v_4846_0;
  wire [2:0] v_4847_0;
  reg [2:0] v_4848_0 = 3'h0;
  wire [0:0] v_4849_0;
  wire [0:0] v_4850_0;
  wire [0:0] v_4851_0;
  wire [2:0] v_4852_0;
  wire [2:0] v_4853_0;
  wire [2:0] v_4854_0;
  reg [2:0] v_4855_0 = 3'h0;
  wire [0:0] v_4856_0;
  wire [0:0] v_4857_0;
  wire [0:0] v_4858_0;
  wire [2:0] v_4859_0;
  wire [2:0] v_4860_0;
  wire [2:0] v_4861_0;
  reg [2:0] v_4862_0 = 3'h0;
  wire [0:0] v_4863_0;
  wire [0:0] v_4864_0;
  wire [0:0] v_4865_0;
  wire [2:0] v_4866_0;
  wire [2:0] v_4867_0;
  wire [2:0] v_4868_0;
  reg [2:0] v_4869_0 = 3'h0;
  wire [0:0] v_4870_0;
  wire [0:0] v_4871_0;
  wire [0:0] v_4872_0;
  wire [2:0] v_4873_0;
  wire [2:0] v_4874_0;
  wire [2:0] v_4875_0;
  reg [2:0] v_4876_0 = 3'h0;
  wire [0:0] v_4877_0;
  wire [0:0] v_4878_0;
  wire [0:0] v_4879_0;
  wire [2:0] v_4880_0;
  wire [2:0] v_4881_0;
  wire [2:0] v_4882_0;
  reg [2:0] v_4883_0 = 3'h0;
  wire [0:0] v_4884_0;
  wire [0:0] v_4885_0;
  wire [0:0] v_4886_0;
  wire [2:0] v_4887_0;
  wire [2:0] v_4888_0;
  wire [2:0] v_4889_0;
  reg [2:0] v_4890_0 = 3'h0;
  wire [0:0] v_4891_0;
  wire [0:0] v_4892_0;
  wire [0:0] v_4893_0;
  wire [2:0] v_4894_0;
  wire [2:0] v_4895_0;
  wire [2:0] v_4896_0;
  reg [2:0] v_4897_0 = 3'h0;
  wire [0:0] v_4898_0;
  wire [0:0] v_4899_0;
  wire [0:0] v_4900_0;
  wire [2:0] v_4901_0;
  wire [2:0] v_4902_0;
  wire [2:0] v_4903_0;
  reg [2:0] v_4904_0 = 3'h0;
  wire [0:0] v_4905_0;
  wire [0:0] v_4906_0;
  wire [0:0] v_4907_0;
  wire [2:0] v_4908_0;
  wire [2:0] v_4909_0;
  wire [2:0] v_4910_0;
  reg [2:0] v_4911_0 = 3'h0;
  wire [0:0] v_4912_0;
  wire [0:0] v_4913_0;
  wire [0:0] v_4914_0;
  wire [2:0] v_4915_0;
  wire [2:0] v_4916_0;
  wire [2:0] v_4917_0;
  reg [2:0] v_4918_0 = 3'h0;
  wire [0:0] v_4919_0;
  wire [0:0] v_4920_0;
  wire [0:0] v_4921_0;
  wire [2:0] v_4922_0;
  wire [2:0] v_4923_0;
  wire [2:0] v_4924_0;
  reg [2:0] v_4925_0 = 3'h0;
  wire [0:0] v_4926_0;
  wire [0:0] v_4927_0;
  wire [0:0] v_4928_0;
  wire [2:0] v_4929_0;
  wire [2:0] v_4930_0;
  wire [2:0] v_4931_0;
  reg [2:0] v_4932_0 = 3'h0;
  wire [0:0] v_4933_0;
  wire [0:0] v_4934_0;
  wire [0:0] v_4935_0;
  wire [2:0] v_4936_0;
  wire [2:0] v_4937_0;
  wire [2:0] v_4938_0;
  reg [2:0] v_4939_0 = 3'h0;
  wire [0:0] v_4940_0;
  wire [0:0] v_4941_0;
  wire [0:0] v_4942_0;
  wire [2:0] v_4943_0;
  wire [2:0] v_4944_0;
  wire [2:0] v_4945_0;
  reg [2:0] v_4946_0 = 3'h0;
  wire [0:0] v_4947_0;
  wire [0:0] v_4948_0;
  wire [0:0] v_4949_0;
  wire [2:0] v_4950_0;
  wire [2:0] v_4951_0;
  wire [2:0] v_4952_0;
  reg [2:0] v_4953_0 = 3'h0;
  wire [0:0] v_4954_0;
  wire [0:0] v_4955_0;
  wire [0:0] v_4956_0;
  wire [2:0] v_4957_0;
  wire [2:0] v_4958_0;
  wire [2:0] v_4959_0;
  reg [2:0] v_4960_0 = 3'h0;
  wire [0:0] v_4961_0;
  wire [0:0] v_4962_0;
  wire [0:0] v_4963_0;
  wire [2:0] v_4964_0;
  wire [2:0] v_4965_0;
  wire [2:0] v_4966_0;
  reg [2:0] v_4967_0 = 3'h0;
  wire [0:0] v_4968_0;
  wire [0:0] v_4969_0;
  wire [0:0] v_4970_0;
  wire [2:0] v_4971_0;
  wire [2:0] v_4972_0;
  wire [2:0] v_4973_0;
  reg [2:0] v_4974_0 = 3'h0;
  wire [0:0] v_4975_0;
  wire [0:0] v_4976_0;
  wire [0:0] v_4977_0;
  wire [2:0] v_4978_0;
  wire [2:0] v_4979_0;
  wire [2:0] v_4980_0;
  reg [2:0] v_4981_0 = 3'h0;
  wire [0:0] v_4982_0;
  wire [0:0] v_4983_0;
  wire [0:0] v_4984_0;
  wire [2:0] v_4985_0;
  wire [2:0] v_4986_0;
  wire [2:0] v_4987_0;
  reg [2:0] v_4988_0 = 3'h0;
  wire [0:0] v_4989_0;
  wire [0:0] v_4990_0;
  wire [0:0] v_4991_0;
  wire [2:0] v_4992_0;
  wire [2:0] v_4993_0;
  wire [2:0] v_4994_0;
  reg [2:0] v_4995_0 = 3'h0;
  wire [0:0] v_4996_0;
  wire [0:0] v_4997_0;
  wire [0:0] v_4998_0;
  wire [2:0] v_4999_0;
  wire [2:0] v_5000_0;
  wire [2:0] v_5001_0;
  reg [2:0] v_5002_0 = 3'h0;
  wire [0:0] v_5003_0;
  wire [0:0] v_5004_0;
  wire [0:0] v_5005_0;
  wire [2:0] v_5006_0;
  wire [2:0] v_5007_0;
  wire [2:0] v_5008_0;
  reg [2:0] v_5009_0 = 3'h0;
  wire [0:0] v_5010_0;
  wire [0:0] v_5011_0;
  wire [0:0] v_5012_0;
  wire [2:0] v_5013_0;
  wire [2:0] v_5014_0;
  wire [2:0] v_5015_0;
  reg [2:0] v_5016_0 = 3'h0;
  wire [0:0] v_5017_0;
  wire [0:0] v_5018_0;
  wire [0:0] v_5019_0;
  wire [2:0] v_5020_0;
  wire [2:0] v_5021_0;
  wire [2:0] v_5022_0;
  reg [2:0] v_5023_0 = 3'h0;
  wire [0:0] v_5024_0;
  wire [0:0] v_5025_0;
  wire [0:0] v_5026_0;
  wire [2:0] v_5027_0;
  wire [2:0] v_5028_0;
  wire [2:0] v_5029_0;
  reg [2:0] v_5030_0 = 3'h0;
  wire [0:0] v_5031_0;
  wire [0:0] v_5032_0;
  wire [0:0] v_5033_0;
  wire [2:0] v_5034_0;
  wire [2:0] v_5035_0;
  wire [2:0] v_5036_0;
  reg [2:0] v_5037_0 = 3'h0;
  wire [0:0] v_5038_0;
  wire [0:0] v_5039_0;
  wire [0:0] v_5040_0;
  wire [2:0] v_5041_0;
  wire [2:0] v_5042_0;
  wire [2:0] v_5043_0;
  reg [2:0] v_5044_0 = 3'h0;
  wire [0:0] v_5045_0;
  wire [0:0] v_5046_0;
  wire [0:0] v_5047_0;
  wire [2:0] v_5048_0;
  wire [2:0] v_5049_0;
  wire [2:0] v_5050_0;
  reg [2:0] v_5051_0 = 3'h0;
  wire [0:0] v_5052_0;
  wire [0:0] v_5053_0;
  wire [0:0] v_5054_0;
  wire [2:0] v_5055_0;
  wire [2:0] v_5056_0;
  wire [2:0] v_5057_0;
  reg [2:0] v_5058_0 = 3'h0;
  wire [0:0] v_5059_0;
  wire [0:0] v_5060_0;
  wire [0:0] v_5061_0;
  wire [2:0] v_5062_0;
  wire [2:0] v_5063_0;
  wire [2:0] v_5064_0;
  reg [2:0] v_5065_0 = 3'h0;
  wire [0:0] v_5066_0;
  wire [0:0] v_5067_0;
  wire [0:0] v_5068_0;
  wire [2:0] v_5069_0;
  wire [2:0] v_5070_0;
  wire [2:0] v_5071_0;
  reg [2:0] v_5072_0 = 3'h0;
  wire [0:0] v_5073_0;
  wire [0:0] v_5074_0;
  wire [0:0] v_5075_0;
  wire [2:0] v_5076_0;
  wire [2:0] v_5077_0;
  wire [2:0] v_5078_0;
  reg [2:0] v_5079_0 = 3'h0;
  wire [0:0] v_5080_0;
  wire [0:0] v_5081_0;
  wire [0:0] v_5082_0;
  wire [2:0] v_5083_0;
  wire [2:0] v_5084_0;
  wire [2:0] v_5085_0;
  reg [2:0] v_5086_0 = 3'h0;
  wire [0:0] v_5087_0;
  wire [0:0] v_5088_0;
  wire [0:0] v_5089_0;
  wire [2:0] v_5090_0;
  wire [2:0] v_5091_0;
  wire [2:0] v_5092_0;
  reg [2:0] v_5093_0 = 3'h0;
  wire [0:0] v_5094_0;
  wire [0:0] v_5095_0;
  wire [0:0] v_5096_0;
  wire [2:0] v_5097_0;
  wire [2:0] v_5098_0;
  wire [2:0] v_5099_0;
  reg [2:0] v_5100_0 = 3'h0;
  wire [0:0] v_5101_0;
  wire [0:0] v_5102_0;
  wire [0:0] v_5103_0;
  wire [2:0] v_5104_0;
  wire [2:0] v_5105_0;
  wire [2:0] v_5106_0;
  reg [2:0] v_5107_0 = 3'h0;
  wire [0:0] v_5108_0;
  wire [0:0] v_5109_0;
  wire [0:0] v_5110_0;
  wire [2:0] v_5111_0;
  wire [2:0] v_5112_0;
  wire [2:0] v_5113_0;
  reg [2:0] v_5114_0 = 3'h0;
  wire [0:0] v_5115_0;
  wire [0:0] v_5116_0;
  wire [0:0] v_5117_0;
  wire [2:0] v_5118_0;
  wire [2:0] v_5119_0;
  wire [2:0] v_5120_0;
  reg [2:0] v_5121_0 = 3'h0;
  wire [0:0] v_5122_0;
  wire [0:0] v_5123_0;
  wire [0:0] v_5124_0;
  wire [2:0] v_5125_0;
  wire [2:0] v_5126_0;
  wire [2:0] v_5127_0;
  reg [2:0] v_5128_0 = 3'h0;
  wire [0:0] v_5129_0;
  wire [0:0] v_5130_0;
  wire [0:0] v_5131_0;
  wire [2:0] v_5132_0;
  wire [2:0] v_5133_0;
  wire [2:0] v_5134_0;
  reg [2:0] v_5135_0 = 3'h0;
  wire [0:0] v_5136_0;
  wire [0:0] v_5137_0;
  wire [0:0] v_5138_0;
  wire [2:0] v_5139_0;
  wire [2:0] v_5140_0;
  wire [2:0] v_5141_0;
  reg [2:0] v_5142_0 = 3'h0;
  wire [0:0] v_5143_0;
  wire [0:0] v_5144_0;
  wire [0:0] v_5145_0;
  wire [2:0] v_5146_0;
  wire [2:0] v_5147_0;
  wire [2:0] v_5148_0;
  reg [2:0] v_5149_0 = 3'h0;
  wire [0:0] v_5150_0;
  wire [0:0] v_5151_0;
  wire [0:0] v_5152_0;
  wire [2:0] v_5153_0;
  wire [2:0] v_5154_0;
  wire [2:0] v_5155_0;
  reg [2:0] v_5156_0 = 3'h0;
  wire [0:0] v_5157_0;
  wire [0:0] v_5158_0;
  wire [0:0] v_5159_0;
  wire [2:0] v_5160_0;
  wire [2:0] v_5161_0;
  wire [2:0] v_5162_0;
  reg [2:0] v_5163_0 = 3'h0;
  wire [0:0] v_5164_0;
  wire [0:0] v_5165_0;
  wire [0:0] v_5166_0;
  wire [2:0] v_5167_0;
  wire [2:0] v_5168_0;
  wire [2:0] v_5169_0;
  reg [2:0] v_5170_0 = 3'h0;
  wire [0:0] v_5171_0;
  wire [0:0] v_5172_0;
  wire [0:0] v_5173_0;
  wire [2:0] v_5174_0;
  wire [2:0] v_5175_0;
  wire [2:0] v_5176_0;
  reg [2:0] v_5177_0 = 3'h0;
  wire [0:0] v_5178_0;
  wire [0:0] v_5179_0;
  wire [0:0] v_5180_0;
  wire [2:0] v_5181_0;
  wire [2:0] v_5182_0;
  wire [2:0] v_5183_0;
  reg [2:0] v_5184_0 = 3'h0;
  wire [0:0] v_5185_0;
  wire [0:0] v_5186_0;
  wire [0:0] v_5187_0;
  wire [2:0] v_5188_0;
  wire [2:0] v_5189_0;
  wire [2:0] v_5190_0;
  reg [2:0] v_5191_0 = 3'h0;
  wire [0:0] v_5192_0;
  wire [0:0] v_5193_0;
  wire [0:0] v_5194_0;
  wire [2:0] v_5195_0;
  wire [2:0] v_5196_0;
  wire [2:0] v_5197_0;
  reg [2:0] v_5198_0 = 3'h0;
  wire [0:0] v_5199_0;
  wire [0:0] v_5200_0;
  wire [0:0] v_5201_0;
  wire [2:0] v_5202_0;
  wire [2:0] v_5203_0;
  wire [2:0] v_5204_0;
  reg [2:0] v_5205_0 = 3'h0;
  wire [0:0] v_5206_0;
  wire [0:0] v_5207_0;
  wire [0:0] v_5208_0;
  wire [2:0] v_5209_0;
  wire [2:0] v_5210_0;
  wire [2:0] v_5211_0;
  reg [2:0] v_5212_0 = 3'h0;
  wire [0:0] v_5213_0;
  wire [0:0] v_5214_0;
  wire [0:0] v_5215_0;
  wire [2:0] v_5216_0;
  wire [2:0] v_5217_0;
  wire [2:0] v_5218_0;
  reg [2:0] v_5219_0 = 3'h0;
  wire [0:0] v_5220_0;
  wire [0:0] v_5221_0;
  wire [0:0] v_5222_0;
  wire [2:0] v_5223_0;
  wire [2:0] v_5224_0;
  wire [2:0] v_5225_0;
  reg [2:0] v_5226_0 = 3'h0;
  wire [0:0] v_5227_0;
  wire [0:0] v_5228_0;
  wire [0:0] v_5229_0;
  wire [2:0] v_5230_0;
  wire [2:0] v_5231_0;
  wire [2:0] v_5232_0;
  reg [2:0] v_5233_0 = 3'h0;
  wire [0:0] v_5234_0;
  wire [0:0] v_5235_0;
  wire [0:0] v_5236_0;
  wire [2:0] v_5237_0;
  wire [2:0] v_5238_0;
  wire [2:0] v_5239_0;
  reg [2:0] v_5240_0 = 3'h0;
  wire [0:0] v_5241_0;
  wire [0:0] v_5242_0;
  wire [0:0] v_5243_0;
  wire [2:0] v_5244_0;
  wire [2:0] v_5245_0;
  wire [2:0] v_5246_0;
  reg [2:0] v_5247_0 = 3'h0;
  wire [0:0] v_5248_0;
  wire [0:0] v_5249_0;
  wire [0:0] v_5250_0;
  wire [2:0] v_5251_0;
  wire [2:0] v_5252_0;
  wire [2:0] v_5253_0;
  reg [2:0] v_5254_0 = 3'h0;
  wire [0:0] v_5255_0;
  wire [0:0] v_5256_0;
  wire [0:0] v_5257_0;
  wire [2:0] v_5258_0;
  wire [2:0] v_5259_0;
  wire [2:0] v_5260_0;
  reg [2:0] v_5261_0 = 3'h0;
  wire [0:0] v_5262_0;
  wire [0:0] v_5263_0;
  wire [0:0] v_5264_0;
  wire [2:0] v_5265_0;
  wire [2:0] v_5266_0;
  wire [2:0] v_5267_0;
  reg [2:0] v_5268_0 = 3'h0;
  wire [0:0] v_5269_0;
  wire [0:0] v_5270_0;
  wire [0:0] v_5271_0;
  wire [2:0] v_5272_0;
  wire [2:0] v_5273_0;
  wire [2:0] v_5274_0;
  reg [2:0] v_5275_0 = 3'h0;
  wire [0:0] v_5276_0;
  wire [0:0] v_5277_0;
  wire [0:0] v_5278_0;
  wire [2:0] v_5279_0;
  wire [2:0] v_5280_0;
  wire [2:0] v_5281_0;
  reg [2:0] v_5282_0 = 3'h0;
  wire [0:0] v_5283_0;
  wire [0:0] v_5284_0;
  wire [0:0] v_5285_0;
  wire [2:0] v_5286_0;
  wire [2:0] v_5287_0;
  wire [2:0] v_5288_0;
  reg [2:0] v_5289_0 = 3'h0;
  wire [0:0] v_5290_0;
  wire [0:0] v_5291_0;
  wire [0:0] v_5292_0;
  wire [2:0] v_5293_0;
  wire [2:0] v_5294_0;
  wire [2:0] v_5295_0;
  reg [2:0] v_5296_0 = 3'h0;
  wire [0:0] v_5297_0;
  wire [0:0] v_5298_0;
  wire [0:0] v_5299_0;
  wire [2:0] v_5300_0;
  wire [2:0] v_5301_0;
  wire [2:0] v_5302_0;
  reg [2:0] v_5303_0 = 3'h0;
  wire [0:0] v_5304_0;
  wire [0:0] v_5305_0;
  wire [0:0] v_5306_0;
  wire [2:0] v_5307_0;
  wire [2:0] v_5308_0;
  wire [2:0] v_5309_0;
  reg [2:0] v_5310_0 = 3'h0;
  wire [0:0] v_5311_0;
  wire [0:0] v_5312_0;
  wire [0:0] v_5313_0;
  wire [2:0] v_5314_0;
  wire [2:0] v_5315_0;
  wire [2:0] v_5316_0;
  reg [2:0] v_5317_0 = 3'h0;
  wire [0:0] v_5318_0;
  wire [0:0] v_5319_0;
  wire [0:0] v_5320_0;
  wire [2:0] v_5321_0;
  wire [2:0] v_5322_0;
  wire [2:0] v_5323_0;
  reg [2:0] v_5324_0 = 3'h0;
  wire [0:0] v_5325_0;
  wire [0:0] v_5326_0;
  wire [0:0] v_5327_0;
  wire [2:0] v_5328_0;
  wire [2:0] v_5329_0;
  wire [2:0] v_5330_0;
  reg [2:0] v_5331_0 = 3'h0;
  wire [0:0] v_5332_0;
  wire [0:0] v_5333_0;
  wire [0:0] v_5334_0;
  wire [2:0] v_5335_0;
  wire [2:0] v_5336_0;
  wire [2:0] v_5337_0;
  reg [2:0] v_5338_0 = 3'h0;
  wire [0:0] v_5339_0;
  wire [0:0] v_5340_0;
  wire [0:0] v_5341_0;
  wire [2:0] v_5342_0;
  wire [2:0] v_5343_0;
  wire [2:0] v_5344_0;
  reg [2:0] v_5345_0 = 3'h0;
  wire [0:0] v_5346_0;
  wire [0:0] v_5347_0;
  wire [0:0] v_5348_0;
  wire [2:0] v_5349_0;
  wire [2:0] v_5350_0;
  wire [2:0] v_5351_0;
  reg [2:0] v_5352_0 = 3'h0;
  wire [0:0] v_5353_0;
  wire [0:0] v_5354_0;
  wire [0:0] v_5355_0;
  wire [2:0] v_5356_0;
  wire [2:0] v_5357_0;
  wire [2:0] v_5358_0;
  reg [2:0] v_5359_0 = 3'h0;
  wire [0:0] v_5360_0;
  wire [0:0] v_5361_0;
  wire [0:0] v_5362_0;
  wire [2:0] v_5363_0;
  wire [2:0] v_5364_0;
  wire [2:0] v_5365_0;
  reg [2:0] v_5366_0 = 3'h0;
  wire [0:0] v_5367_0;
  wire [0:0] v_5368_0;
  wire [0:0] v_5369_0;
  wire [2:0] v_5370_0;
  wire [2:0] v_5371_0;
  wire [2:0] v_5372_0;
  reg [2:0] v_5373_0 = 3'h0;
  wire [0:0] v_5374_0;
  wire [0:0] v_5375_0;
  wire [0:0] v_5376_0;
  wire [2:0] v_5377_0;
  wire [2:0] v_5378_0;
  wire [2:0] v_5379_0;
  reg [2:0] v_5380_0 = 3'h0;
  wire [0:0] v_5381_0;
  wire [0:0] v_5382_0;
  wire [0:0] v_5383_0;
  wire [2:0] v_5384_0;
  wire [2:0] v_5385_0;
  wire [2:0] v_5386_0;
  reg [2:0] v_5387_0 = 3'h0;
  wire [0:0] v_5388_0;
  wire [0:0] v_5389_0;
  wire [0:0] v_5390_0;
  wire [2:0] v_5391_0;
  wire [2:0] v_5392_0;
  wire [2:0] v_5393_0;
  reg [2:0] v_5394_0 = 3'h0;
  wire [0:0] v_5395_0;
  wire [0:0] v_5396_0;
  wire [0:0] v_5397_0;
  wire [2:0] v_5398_0;
  wire [2:0] v_5399_0;
  wire [2:0] v_5400_0;
  reg [2:0] v_5401_0 = 3'h0;
  wire [0:0] v_5402_0;
  wire [0:0] v_5403_0;
  wire [0:0] v_5404_0;
  wire [2:0] v_5405_0;
  wire [2:0] v_5406_0;
  wire [2:0] v_5407_0;
  reg [2:0] v_5408_0 = 3'h0;
  wire [0:0] v_5409_0;
  wire [0:0] v_5410_0;
  wire [0:0] v_5411_0;
  wire [2:0] v_5412_0;
  wire [2:0] v_5413_0;
  wire [2:0] v_5414_0;
  reg [2:0] v_5415_0 = 3'h0;
  wire [0:0] v_5416_0;
  wire [0:0] v_5417_0;
  wire [0:0] v_5418_0;
  wire [2:0] v_5419_0;
  wire [2:0] v_5420_0;
  wire [2:0] v_5421_0;
  reg [2:0] v_5422_0 = 3'h0;
  wire [0:0] v_5423_0;
  wire [0:0] v_5424_0;
  wire [0:0] v_5425_0;
  wire [2:0] v_5426_0;
  wire [2:0] v_5427_0;
  wire [2:0] v_5428_0;
  reg [2:0] v_5429_0 = 3'h0;
  wire [0:0] v_5430_0;
  wire [0:0] v_5431_0;
  wire [0:0] v_5432_0;
  wire [2:0] v_5433_0;
  wire [2:0] v_5434_0;
  wire [2:0] v_5435_0;
  reg [2:0] v_5436_0 = 3'h0;
  wire [0:0] v_5437_0;
  wire [0:0] v_5438_0;
  wire [0:0] v_5439_0;
  wire [2:0] v_5440_0;
  wire [2:0] v_5441_0;
  wire [2:0] v_5442_0;
  reg [2:0] v_5443_0 = 3'h0;
  wire [0:0] v_5444_0;
  wire [0:0] v_5445_0;
  wire [0:0] v_5446_0;
  wire [2:0] v_5447_0;
  wire [2:0] v_5448_0;
  wire [2:0] v_5449_0;
  reg [2:0] v_5450_0 = 3'h0;
  wire [0:0] v_5451_0;
  wire [0:0] v_5452_0;
  wire [0:0] v_5453_0;
  wire [2:0] v_5454_0;
  wire [2:0] v_5455_0;
  wire [2:0] v_5456_0;
  reg [2:0] v_5457_0 = 3'h0;
  wire [0:0] v_5458_0;
  wire [0:0] v_5459_0;
  wire [0:0] v_5460_0;
  wire [2:0] v_5461_0;
  wire [2:0] v_5462_0;
  wire [2:0] v_5463_0;
  reg [2:0] v_5464_0 = 3'h0;
  wire [0:0] v_5465_0;
  wire [0:0] v_5466_0;
  wire [0:0] v_5467_0;
  wire [2:0] v_5468_0;
  wire [2:0] v_5469_0;
  wire [2:0] v_5470_0;
  reg [2:0] v_5471_0 = 3'h0;
  wire [0:0] v_5472_0;
  wire [0:0] v_5473_0;
  wire [0:0] v_5474_0;
  wire [2:0] v_5475_0;
  wire [2:0] v_5476_0;
  wire [2:0] v_5477_0;
  reg [2:0] v_5478_0 = 3'h0;
  wire [0:0] v_5479_0;
  wire [0:0] v_5480_0;
  wire [0:0] v_5481_0;
  wire [2:0] v_5482_0;
  wire [2:0] v_5483_0;
  wire [2:0] v_5484_0;
  reg [2:0] v_5485_0 = 3'h0;
  wire [0:0] v_5486_0;
  wire [0:0] v_5487_0;
  wire [0:0] v_5488_0;
  wire [2:0] v_5489_0;
  wire [2:0] v_5490_0;
  wire [2:0] v_5491_0;
  reg [2:0] v_5492_0 = 3'h0;
  wire [0:0] v_5493_0;
  wire [0:0] v_5494_0;
  wire [0:0] v_5495_0;
  wire [2:0] v_5496_0;
  wire [2:0] v_5497_0;
  wire [2:0] v_5498_0;
  reg [2:0] v_5499_0 = 3'h0;
  wire [0:0] v_5500_0;
  wire [0:0] v_5501_0;
  wire [0:0] v_5502_0;
  wire [2:0] v_5503_0;
  wire [2:0] v_5504_0;
  wire [2:0] v_5505_0;
  reg [2:0] v_5506_0 = 3'h0;
  wire [0:0] v_5507_0;
  wire [0:0] v_5508_0;
  wire [0:0] v_5509_0;
  wire [2:0] v_5510_0;
  wire [2:0] v_5511_0;
  wire [2:0] v_5512_0;
  reg [2:0] v_5513_0 = 3'h0;
  wire [0:0] v_5514_0;
  wire [0:0] v_5515_0;
  wire [0:0] v_5516_0;
  wire [2:0] v_5517_0;
  wire [2:0] v_5518_0;
  wire [2:0] v_5519_0;
  reg [2:0] v_5520_0 = 3'h0;
  wire [0:0] v_5521_0;
  wire [0:0] v_5522_0;
  wire [0:0] v_5523_0;
  wire [2:0] v_5524_0;
  wire [2:0] v_5525_0;
  wire [2:0] v_5526_0;
  reg [2:0] v_5527_0 = 3'h0;
  wire [0:0] v_5528_0;
  wire [0:0] v_5529_0;
  wire [0:0] v_5530_0;
  wire [2:0] v_5531_0;
  wire [2:0] v_5532_0;
  wire [2:0] v_5533_0;
  reg [2:0] v_5534_0 = 3'h0;
  wire [0:0] v_5535_0;
  wire [0:0] v_5536_0;
  wire [0:0] v_5537_0;
  wire [2:0] v_5538_0;
  wire [2:0] v_5539_0;
  wire [2:0] v_5540_0;
  reg [2:0] v_5541_0 = 3'h0;
  wire [0:0] v_5542_0;
  wire [0:0] v_5543_0;
  wire [0:0] v_5544_0;
  wire [2:0] v_5545_0;
  wire [2:0] v_5546_0;
  wire [2:0] v_5547_0;
  reg [2:0] v_5548_0 = 3'h0;
  wire [0:0] v_5549_0;
  wire [0:0] v_5550_0;
  wire [0:0] v_5551_0;
  wire [2:0] v_5552_0;
  wire [2:0] v_5553_0;
  wire [2:0] v_5554_0;
  reg [2:0] v_5555_0 = 3'h0;
  wire [0:0] v_5556_0;
  wire [0:0] v_5557_0;
  wire [0:0] v_5558_0;
  wire [2:0] v_5559_0;
  wire [2:0] v_5560_0;
  wire [2:0] v_5561_0;
  reg [2:0] v_5562_0 = 3'h0;
  wire [0:0] v_5563_0;
  wire [0:0] v_5564_0;
  wire [0:0] v_5565_0;
  wire [2:0] v_5566_0;
  wire [2:0] v_5567_0;
  wire [2:0] v_5568_0;
  reg [2:0] v_5569_0 = 3'h0;
  wire [0:0] v_5570_0;
  wire [0:0] v_5571_0;
  wire [0:0] v_5572_0;
  wire [2:0] v_5573_0;
  wire [2:0] v_5574_0;
  wire [2:0] v_5575_0;
  reg [2:0] v_5576_0 = 3'h0;
  wire [0:0] v_5577_0;
  wire [0:0] v_5578_0;
  wire [0:0] v_5579_0;
  wire [2:0] v_5580_0;
  wire [2:0] v_5581_0;
  wire [2:0] v_5582_0;
  reg [2:0] v_5583_0 = 3'h0;
  wire [0:0] v_5584_0;
  wire [0:0] v_5585_0;
  wire [0:0] v_5586_0;
  wire [2:0] v_5587_0;
  wire [2:0] v_5588_0;
  wire [2:0] v_5589_0;
  reg [2:0] v_5590_0 = 3'h0;
  wire [0:0] v_5591_0;
  wire [0:0] v_5592_0;
  wire [0:0] v_5593_0;
  wire [2:0] v_5594_0;
  wire [2:0] v_5595_0;
  wire [2:0] v_5596_0;
  reg [2:0] v_5597_0 = 3'h0;
  wire [0:0] v_5598_0;
  wire [0:0] v_5599_0;
  wire [0:0] v_5600_0;
  wire [2:0] v_5601_0;
  wire [2:0] v_5602_0;
  wire [2:0] v_5603_0;
  reg [2:0] v_5604_0 = 3'h0;
  wire [0:0] v_5605_0;
  wire [0:0] v_5606_0;
  wire [0:0] v_5607_0;
  wire [2:0] v_5608_0;
  wire [2:0] v_5609_0;
  wire [2:0] v_5610_0;
  reg [2:0] v_5611_0 = 3'h0;
  wire [0:0] v_5612_0;
  wire [0:0] v_5613_0;
  wire [0:0] v_5614_0;
  wire [2:0] v_5615_0;
  wire [2:0] v_5616_0;
  wire [2:0] v_5617_0;
  reg [2:0] v_5618_0 = 3'h0;
  wire [0:0] v_5619_0;
  wire [0:0] v_5620_0;
  wire [0:0] v_5621_0;
  wire [2:0] v_5622_0;
  wire [2:0] v_5623_0;
  wire [2:0] v_5624_0;
  reg [2:0] v_5625_0 = 3'h0;
  wire [0:0] v_5626_0;
  wire [0:0] v_5627_0;
  wire [0:0] v_5628_0;
  wire [2:0] v_5629_0;
  wire [2:0] v_5630_0;
  wire [2:0] v_5631_0;
  reg [2:0] v_5632_0 = 3'h0;
  wire [0:0] v_5633_0;
  wire [0:0] v_5634_0;
  wire [0:0] v_5635_0;
  wire [2:0] v_5636_0;
  wire [2:0] v_5637_0;
  wire [2:0] v_5638_0;
  reg [2:0] v_5639_0 = 3'h0;
  wire [0:0] v_5640_0;
  wire [0:0] v_5641_0;
  wire [0:0] v_5642_0;
  wire [2:0] v_5643_0;
  wire [2:0] v_5644_0;
  wire [2:0] v_5645_0;
  reg [2:0] v_5646_0 = 3'h0;
  wire [0:0] v_5647_0;
  wire [0:0] v_5648_0;
  wire [0:0] v_5649_0;
  wire [2:0] v_5650_0;
  wire [2:0] v_5651_0;
  wire [2:0] v_5652_0;
  reg [2:0] v_5653_0 = 3'h0;
  wire [0:0] v_5654_0;
  wire [0:0] v_5655_0;
  wire [0:0] v_5656_0;
  wire [2:0] v_5657_0;
  wire [2:0] v_5658_0;
  wire [2:0] v_5659_0;
  reg [2:0] v_5660_0 = 3'h0;
  wire [0:0] v_5661_0;
  wire [0:0] v_5662_0;
  wire [0:0] v_5663_0;
  wire [2:0] v_5664_0;
  wire [2:0] v_5665_0;
  wire [2:0] v_5666_0;
  reg [2:0] v_5667_0 = 3'h0;
  wire [0:0] v_5668_0;
  wire [0:0] v_5669_0;
  wire [0:0] v_5670_0;
  wire [2:0] v_5671_0;
  wire [2:0] v_5672_0;
  wire [2:0] v_5673_0;
  reg [2:0] v_5674_0 = 3'h0;
  wire [0:0] v_5675_0;
  wire [0:0] v_5676_0;
  wire [0:0] v_5677_0;
  wire [2:0] v_5678_0;
  wire [2:0] v_5679_0;
  wire [2:0] v_5680_0;
  reg [2:0] v_5681_0 = 3'h0;
  wire [0:0] v_5682_0;
  wire [0:0] v_5683_0;
  wire [0:0] v_5684_0;
  wire [2:0] v_5685_0;
  wire [2:0] v_5686_0;
  wire [2:0] v_5687_0;
  reg [2:0] v_5688_0 = 3'h0;
  wire [0:0] v_5689_0;
  wire [0:0] v_5690_0;
  wire [0:0] v_5691_0;
  wire [2:0] v_5692_0;
  wire [2:0] v_5693_0;
  wire [2:0] v_5694_0;
  reg [2:0] v_5695_0 = 3'h0;
  wire [0:0] v_5696_0;
  wire [0:0] v_5697_0;
  wire [0:0] v_5698_0;
  wire [2:0] v_5699_0;
  wire [2:0] v_5700_0;
  wire [2:0] v_5701_0;
  reg [2:0] v_5702_0 = 3'h0;
  wire [0:0] v_5703_0;
  wire [0:0] v_5704_0;
  wire [0:0] v_5705_0;
  wire [2:0] v_5706_0;
  wire [2:0] v_5707_0;
  wire [2:0] v_5708_0;
  reg [2:0] v_5709_0 = 3'h0;
  wire [0:0] v_5710_0;
  wire [0:0] v_5711_0;
  wire [0:0] v_5712_0;
  wire [2:0] v_5713_0;
  wire [2:0] v_5714_0;
  wire [2:0] v_5715_0;
  reg [2:0] v_5716_0 = 3'h0;
  wire [0:0] v_5717_0;
  wire [0:0] v_5718_0;
  wire [0:0] v_5719_0;
  wire [2:0] v_5720_0;
  wire [2:0] v_5721_0;
  wire [2:0] v_5722_0;
  reg [2:0] v_5723_0 = 3'h0;
  wire [0:0] v_5724_0;
  wire [0:0] v_5725_0;
  wire [0:0] v_5726_0;
  wire [2:0] v_5727_0;
  wire [2:0] v_5728_0;
  wire [2:0] v_5729_0;
  reg [2:0] v_5730_0 = 3'h0;
  wire [0:0] v_5731_0;
  wire [0:0] v_5732_0;
  wire [0:0] v_5733_0;
  wire [2:0] v_5734_0;
  wire [2:0] v_5735_0;
  wire [2:0] v_5736_0;
  reg [2:0] v_5737_0 = 3'h0;
  wire [0:0] v_5738_0;
  wire [0:0] v_5739_0;
  wire [0:0] v_5740_0;
  wire [2:0] v_5741_0;
  wire [2:0] v_5742_0;
  wire [2:0] v_5743_0;
  reg [2:0] v_5744_0 = 3'h0;
  wire [0:0] v_5745_0;
  wire [0:0] v_5746_0;
  wire [0:0] v_5747_0;
  wire [2:0] v_5748_0;
  wire [2:0] v_5749_0;
  wire [2:0] v_5750_0;
  reg [2:0] v_5751_0 = 3'h0;
  wire [0:0] v_5752_0;
  wire [0:0] v_5753_0;
  wire [0:0] v_5754_0;
  wire [2:0] v_5755_0;
  wire [2:0] v_5756_0;
  wire [2:0] v_5757_0;
  reg [2:0] v_5758_0 = 3'h0;
  wire [0:0] v_5759_0;
  wire [0:0] v_5760_0;
  wire [0:0] v_5761_0;
  wire [2:0] v_5762_0;
  wire [2:0] v_5763_0;
  wire [2:0] v_5764_0;
  reg [2:0] v_5765_0 = 3'h0;
  wire [0:0] v_5766_0;
  wire [0:0] v_5767_0;
  wire [0:0] v_5768_0;
  wire [2:0] v_5769_0;
  wire [2:0] v_5770_0;
  wire [2:0] v_5771_0;
  reg [2:0] v_5772_0 = 3'h0;
  wire [0:0] v_5773_0;
  wire [0:0] v_5774_0;
  wire [0:0] v_5775_0;
  wire [2:0] v_5776_0;
  wire [2:0] v_5777_0;
  wire [2:0] v_5778_0;
  reg [2:0] v_5779_0 = 3'h0;
  wire [0:0] v_5780_0;
  wire [0:0] v_5781_0;
  wire [0:0] v_5782_0;
  wire [2:0] v_5783_0;
  wire [2:0] v_5784_0;
  wire [2:0] v_5785_0;
  reg [2:0] v_5786_0 = 3'h0;
  wire [0:0] v_5787_0;
  wire [0:0] v_5788_0;
  wire [0:0] v_5789_0;
  wire [2:0] v_5790_0;
  wire [2:0] v_5791_0;
  wire [2:0] v_5792_0;
  reg [2:0] v_5793_0 = 3'h0;
  wire [0:0] v_5794_0;
  wire [0:0] v_5795_0;
  wire [0:0] v_5796_0;
  wire [2:0] v_5797_0;
  wire [2:0] v_5798_0;
  wire [2:0] v_5799_0;
  reg [2:0] v_5800_0 = 3'h0;
  wire [0:0] v_5801_0;
  wire [0:0] v_5802_0;
  wire [0:0] v_5803_0;
  wire [2:0] v_5804_0;
  wire [2:0] v_5805_0;
  wire [2:0] v_5806_0;
  reg [2:0] v_5807_0 = 3'h0;
  wire [0:0] v_5808_0;
  wire [0:0] v_5809_0;
  wire [0:0] v_5810_0;
  wire [2:0] v_5811_0;
  wire [2:0] v_5812_0;
  wire [2:0] v_5813_0;
  reg [2:0] v_5814_0 = 3'h0;
  wire [0:0] v_5815_0;
  wire [0:0] v_5816_0;
  wire [0:0] v_5817_0;
  wire [2:0] v_5818_0;
  wire [2:0] v_5819_0;
  wire [2:0] v_5820_0;
  reg [2:0] v_5821_0 = 3'h0;
  wire [0:0] v_5822_0;
  wire [0:0] v_5823_0;
  wire [0:0] v_5824_0;
  wire [2:0] v_5825_0;
  wire [2:0] v_5826_0;
  wire [2:0] v_5827_0;
  reg [2:0] v_5828_0 = 3'h0;
  wire [0:0] v_5829_0;
  wire [0:0] v_5830_0;
  wire [0:0] v_5831_0;
  wire [2:0] v_5832_0;
  wire [2:0] v_5833_0;
  wire [2:0] v_5834_0;
  reg [2:0] v_5835_0 = 3'h0;
  wire [0:0] v_5836_0;
  wire [0:0] v_5837_0;
  wire [0:0] v_5838_0;
  wire [2:0] v_5839_0;
  wire [2:0] v_5840_0;
  wire [2:0] v_5841_0;
  reg [2:0] v_5842_0 = 3'h0;
  wire [0:0] v_5843_0;
  wire [0:0] v_5844_0;
  wire [0:0] v_5845_0;
  wire [2:0] v_5846_0;
  wire [2:0] v_5847_0;
  wire [2:0] v_5848_0;
  reg [2:0] v_5849_0 = 3'h0;
  wire [0:0] v_5850_0;
  wire [0:0] v_5851_0;
  wire [0:0] v_5852_0;
  wire [2:0] v_5853_0;
  wire [2:0] v_5854_0;
  wire [2:0] v_5855_0;
  reg [2:0] v_5856_0 = 3'h0;
  wire [0:0] v_5857_0;
  wire [0:0] v_5858_0;
  wire [0:0] v_5859_0;
  wire [2:0] v_5860_0;
  wire [2:0] v_5861_0;
  wire [2:0] v_5862_0;
  reg [2:0] v_5863_0 = 3'h0;
  wire [0:0] v_5864_0;
  wire [0:0] v_5865_0;
  wire [0:0] v_5866_0;
  wire [2:0] v_5867_0;
  wire [2:0] v_5868_0;
  wire [2:0] v_5869_0;
  reg [2:0] v_5870_0 = 3'h0;
  wire [0:0] v_5871_0;
  wire [0:0] v_5872_0;
  wire [0:0] v_5873_0;
  wire [2:0] v_5874_0;
  wire [2:0] v_5875_0;
  wire [2:0] v_5876_0;
  reg [2:0] v_5877_0 = 3'h0;
  wire [0:0] v_5878_0;
  wire [0:0] v_5879_0;
  wire [0:0] v_5880_0;
  wire [2:0] v_5881_0;
  wire [2:0] v_5882_0;
  wire [2:0] v_5883_0;
  reg [2:0] v_5884_0 = 3'h0;
  wire [0:0] v_5885_0;
  wire [0:0] v_5886_0;
  wire [0:0] v_5887_0;
  wire [2:0] v_5888_0;
  wire [2:0] v_5889_0;
  wire [2:0] v_5890_0;
  reg [2:0] v_5891_0 = 3'h0;
  wire [0:0] v_5892_0;
  wire [0:0] v_5893_0;
  wire [0:0] v_5894_0;
  wire [2:0] v_5895_0;
  wire [2:0] v_5896_0;
  wire [2:0] v_5897_0;
  reg [2:0] v_5898_0 = 3'h0;
  wire [0:0] v_5899_0;
  wire [0:0] v_5900_0;
  wire [0:0] v_5901_0;
  wire [2:0] v_5902_0;
  wire [2:0] v_5903_0;
  wire [2:0] v_5904_0;
  reg [2:0] v_5905_0 = 3'h0;
  wire [0:0] v_5906_0;
  wire [0:0] v_5907_0;
  wire [0:0] v_5908_0;
  wire [2:0] v_5909_0;
  wire [2:0] v_5910_0;
  wire [2:0] v_5911_0;
  reg [2:0] v_5912_0 = 3'h0;
  wire [0:0] v_5913_0;
  wire [0:0] v_5914_0;
  wire [0:0] v_5915_0;
  wire [2:0] v_5916_0;
  wire [2:0] v_5917_0;
  wire [2:0] v_5918_0;
  reg [2:0] v_5919_0 = 3'h0;
  wire [0:0] v_5920_0;
  wire [0:0] v_5921_0;
  wire [0:0] v_5922_0;
  wire [2:0] v_5923_0;
  wire [2:0] v_5924_0;
  wire [2:0] v_5925_0;
  reg [2:0] v_5926_0 = 3'h0;
  wire [0:0] v_5927_0;
  wire [0:0] v_5928_0;
  wire [0:0] v_5929_0;
  wire [2:0] v_5930_0;
  wire [2:0] v_5931_0;
  wire [2:0] v_5932_0;
  reg [2:0] v_5933_0 = 3'h0;
  wire [0:0] v_5934_0;
  wire [0:0] v_5935_0;
  wire [0:0] v_5936_0;
  wire [2:0] v_5937_0;
  wire [2:0] v_5938_0;
  wire [2:0] v_5939_0;
  reg [2:0] v_5940_0 = 3'h0;
  wire [0:0] v_5941_0;
  wire [0:0] v_5942_0;
  wire [0:0] v_5943_0;
  wire [2:0] v_5944_0;
  wire [2:0] v_5945_0;
  wire [2:0] v_5946_0;
  reg [2:0] v_5947_0 = 3'h0;
  wire [0:0] v_5948_0;
  wire [0:0] v_5949_0;
  wire [0:0] v_5950_0;
  wire [2:0] v_5951_0;
  wire [2:0] v_5952_0;
  wire [2:0] v_5953_0;
  reg [2:0] v_5954_0 = 3'h0;
  wire [0:0] v_5955_0;
  wire [0:0] v_5956_0;
  wire [0:0] v_5957_0;
  wire [2:0] v_5958_0;
  wire [2:0] v_5959_0;
  wire [2:0] v_5960_0;
  reg [2:0] v_5961_0 = 3'h0;
  wire [0:0] v_5962_0;
  wire [0:0] v_5963_0;
  wire [0:0] v_5964_0;
  wire [2:0] v_5965_0;
  wire [2:0] v_5966_0;
  wire [2:0] v_5967_0;
  reg [2:0] v_5968_0 = 3'h0;
  wire [0:0] v_5969_0;
  wire [0:0] v_5970_0;
  wire [0:0] v_5971_0;
  wire [2:0] v_5972_0;
  wire [2:0] v_5973_0;
  wire [2:0] v_5974_0;
  reg [2:0] v_5975_0 = 3'h0;
  wire [0:0] v_5976_0;
  wire [0:0] v_5977_0;
  wire [0:0] v_5978_0;
  wire [2:0] v_5979_0;
  wire [2:0] v_5980_0;
  wire [2:0] v_5981_0;
  reg [2:0] v_5982_0 = 3'h0;
  wire [0:0] v_5983_0;
  wire [0:0] v_5984_0;
  wire [0:0] v_5985_0;
  wire [2:0] v_5986_0;
  wire [2:0] v_5987_0;
  wire [2:0] v_5988_0;
  reg [2:0] v_5989_0 = 3'h0;
  wire [0:0] v_5990_0;
  wire [0:0] v_5991_0;
  wire [0:0] v_5992_0;
  wire [2:0] v_5993_0;
  wire [2:0] v_5994_0;
  wire [2:0] v_5995_0;
  reg [2:0] v_5996_0 = 3'h0;
  wire [0:0] v_5997_0;
  wire [0:0] v_5998_0;
  wire [0:0] v_5999_0;
  wire [2:0] v_6000_0;
  wire [2:0] v_6001_0;
  wire [2:0] v_6002_0;
  reg [2:0] v_6003_0 = 3'h0;
  wire [0:0] v_6004_0;
  wire [0:0] v_6005_0;
  wire [0:0] v_6006_0;
  wire [2:0] v_6007_0;
  wire [2:0] v_6008_0;
  wire [2:0] v_6009_0;
  reg [2:0] v_6010_0 = 3'h0;
  wire [0:0] v_6011_0;
  wire [0:0] v_6012_0;
  wire [0:0] v_6013_0;
  wire [2:0] v_6014_0;
  wire [2:0] v_6015_0;
  wire [2:0] v_6016_0;
  reg [2:0] v_6017_0 = 3'h0;
  wire [0:0] v_6018_0;
  wire [0:0] v_6019_0;
  wire [0:0] v_6020_0;
  wire [2:0] v_6021_0;
  wire [2:0] v_6022_0;
  wire [2:0] v_6023_0;
  reg [2:0] v_6024_0 = 3'h0;
  wire [0:0] v_6025_0;
  wire [0:0] v_6026_0;
  wire [0:0] v_6027_0;
  wire [2:0] v_6028_0;
  wire [2:0] v_6029_0;
  wire [2:0] v_6030_0;
  reg [2:0] v_6031_0 = 3'h0;
  wire [0:0] v_6032_0;
  wire [0:0] v_6033_0;
  wire [0:0] v_6034_0;
  wire [2:0] v_6035_0;
  wire [2:0] v_6036_0;
  wire [2:0] v_6037_0;
  reg [2:0] v_6038_0 = 3'h0;
  wire [0:0] v_6039_0;
  wire [0:0] v_6040_0;
  wire [0:0] v_6041_0;
  wire [2:0] v_6042_0;
  wire [2:0] v_6043_0;
  wire [2:0] v_6044_0;
  reg [2:0] v_6045_0 = 3'h0;
  wire [0:0] v_6046_0;
  wire [0:0] v_6047_0;
  wire [0:0] v_6048_0;
  wire [2:0] v_6049_0;
  wire [2:0] v_6050_0;
  wire [2:0] v_6051_0;
  reg [2:0] v_6052_0 = 3'h0;
  wire [0:0] v_6053_0;
  wire [0:0] v_6054_0;
  wire [0:0] v_6055_0;
  wire [2:0] v_6056_0;
  wire [2:0] v_6057_0;
  wire [2:0] v_6058_0;
  reg [2:0] v_6059_0 = 3'h0;
  wire [0:0] v_6060_0;
  wire [0:0] v_6061_0;
  wire [0:0] v_6062_0;
  wire [2:0] v_6063_0;
  wire [2:0] v_6064_0;
  wire [2:0] v_6065_0;
  reg [2:0] v_6066_0 = 3'h0;
  wire [0:0] v_6067_0;
  wire [0:0] v_6068_0;
  wire [0:0] v_6069_0;
  wire [2:0] v_6070_0;
  wire [2:0] v_6071_0;
  wire [2:0] v_6072_0;
  reg [2:0] v_6073_0 = 3'h0;
  wire [0:0] v_6074_0;
  wire [0:0] v_6075_0;
  wire [0:0] v_6076_0;
  wire [2:0] v_6077_0;
  wire [2:0] v_6078_0;
  wire [2:0] v_6079_0;
  reg [2:0] v_6080_0 = 3'h0;
  wire [0:0] v_6081_0;
  wire [0:0] v_6082_0;
  wire [0:0] v_6083_0;
  wire [2:0] v_6084_0;
  wire [2:0] v_6085_0;
  wire [2:0] v_6086_0;
  reg [2:0] v_6087_0 = 3'h0;
  wire [0:0] v_6088_0;
  wire [0:0] v_6089_0;
  wire [0:0] v_6090_0;
  wire [2:0] v_6091_0;
  wire [2:0] v_6092_0;
  wire [2:0] v_6093_0;
  reg [2:0] v_6094_0 = 3'h0;
  wire [0:0] v_6095_0;
  wire [0:0] v_6096_0;
  wire [0:0] v_6097_0;
  wire [2:0] v_6098_0;
  wire [2:0] v_6099_0;
  wire [2:0] v_6100_0;
  reg [2:0] v_6101_0 = 3'h0;
  wire [0:0] v_6102_0;
  wire [0:0] v_6103_0;
  wire [0:0] v_6104_0;
  wire [2:0] v_6105_0;
  wire [2:0] v_6106_0;
  wire [2:0] v_6107_0;
  reg [2:0] v_6108_0 = 3'h0;
  wire [0:0] v_6109_0;
  wire [0:0] v_6110_0;
  wire [0:0] v_6111_0;
  wire [2:0] v_6112_0;
  wire [2:0] v_6113_0;
  wire [2:0] v_6114_0;
  reg [2:0] v_6115_0 = 3'h0;
  wire [0:0] v_6116_0;
  wire [0:0] v_6117_0;
  wire [0:0] v_6118_0;
  wire [2:0] v_6119_0;
  wire [2:0] v_6120_0;
  wire [2:0] v_6121_0;
  reg [2:0] v_6122_0 = 3'h0;
  wire [0:0] v_6123_0;
  wire [0:0] v_6124_0;
  wire [0:0] v_6125_0;
  wire [2:0] v_6126_0;
  wire [2:0] v_6127_0;
  wire [2:0] v_6128_0;
  reg [2:0] v_6129_0 = 3'h0;
  wire [0:0] v_6130_0;
  wire [0:0] v_6131_0;
  wire [0:0] v_6132_0;
  wire [2:0] v_6133_0;
  wire [2:0] v_6134_0;
  wire [2:0] v_6135_0;
  reg [2:0] v_6136_0 = 3'h0;
  wire [0:0] v_6137_0;
  wire [0:0] v_6138_0;
  wire [0:0] v_6139_0;
  wire [2:0] v_6140_0;
  wire [2:0] v_6141_0;
  wire [2:0] v_6142_0;
  reg [2:0] v_6143_0 = 3'h0;
  wire [0:0] v_6144_0;
  wire [0:0] v_6145_0;
  wire [0:0] v_6146_0;
  wire [2:0] v_6147_0;
  wire [2:0] v_6148_0;
  wire [2:0] v_6149_0;
  reg [2:0] v_6150_0 = 3'h0;
  wire [0:0] v_6151_0;
  wire [0:0] v_6152_0;
  wire [0:0] v_6153_0;
  wire [2:0] v_6154_0;
  wire [2:0] v_6155_0;
  wire [2:0] v_6156_0;
  reg [2:0] v_6157_0 = 3'h0;
  wire [0:0] v_6158_0;
  wire [0:0] v_6159_0;
  wire [0:0] v_6160_0;
  wire [2:0] v_6161_0;
  wire [2:0] v_6162_0;
  wire [2:0] v_6163_0;
  reg [2:0] v_6164_0 = 3'h0;
  wire [0:0] v_6165_0;
  wire [0:0] v_6166_0;
  wire [0:0] v_6167_0;
  wire [2:0] v_6168_0;
  wire [2:0] v_6169_0;
  wire [2:0] v_6170_0;
  reg [2:0] v_6171_0 = 3'h0;
  wire [0:0] v_6172_0;
  wire [0:0] v_6173_0;
  wire [0:0] v_6174_0;
  wire [2:0] v_6175_0;
  wire [2:0] v_6176_0;
  wire [2:0] v_6177_0;
  reg [2:0] v_6178_0 = 3'h0;
  wire [0:0] v_6179_0;
  wire [0:0] v_6180_0;
  wire [0:0] v_6181_0;
  wire [2:0] v_6182_0;
  wire [2:0] v_6183_0;
  wire [2:0] v_6184_0;
  reg [2:0] v_6185_0 = 3'h0;
  wire [0:0] v_6186_0;
  wire [0:0] v_6187_0;
  wire [0:0] v_6188_0;
  wire [2:0] v_6189_0;
  wire [2:0] v_6190_0;
  wire [2:0] v_6191_0;
  reg [2:0] v_6192_0 = 3'h0;
  wire [0:0] v_6193_0;
  wire [0:0] v_6194_0;
  wire [0:0] v_6195_0;
  wire [2:0] v_6196_0;
  wire [2:0] v_6197_0;
  wire [2:0] v_6198_0;
  reg [2:0] v_6199_0 = 3'h0;
  wire [0:0] v_6200_0;
  wire [0:0] v_6201_0;
  wire [0:0] v_6202_0;
  wire [2:0] v_6203_0;
  wire [2:0] v_6204_0;
  wire [2:0] v_6205_0;
  reg [2:0] v_6206_0 = 3'h0;
  wire [0:0] v_6207_0;
  wire [0:0] v_6208_0;
  wire [0:0] v_6209_0;
  wire [2:0] v_6210_0;
  wire [2:0] v_6211_0;
  wire [2:0] v_6212_0;
  reg [2:0] v_6213_0 = 3'h0;
  wire [0:0] v_6214_0;
  wire [0:0] v_6215_0;
  wire [0:0] v_6216_0;
  wire [2:0] v_6217_0;
  wire [2:0] v_6218_0;
  wire [2:0] v_6219_0;
  reg [2:0] v_6220_0 = 3'h0;
  wire [0:0] v_6221_0;
  wire [0:0] v_6222_0;
  wire [0:0] v_6223_0;
  wire [2:0] v_6224_0;
  wire [2:0] v_6225_0;
  wire [2:0] v_6226_0;
  reg [2:0] v_6227_0 = 3'h0;
  wire [0:0] v_6228_0;
  wire [0:0] v_6229_0;
  wire [0:0] v_6230_0;
  wire [2:0] v_6231_0;
  wire [2:0] v_6232_0;
  wire [2:0] v_6233_0;
  reg [2:0] v_6234_0 = 3'h0;
  wire [0:0] v_6235_0;
  wire [0:0] v_6236_0;
  wire [0:0] v_6237_0;
  wire [2:0] v_6238_0;
  wire [2:0] v_6239_0;
  wire [2:0] v_6240_0;
  reg [2:0] v_6241_0 = 3'h0;
  wire [0:0] v_6242_0;
  wire [0:0] v_6243_0;
  wire [0:0] v_6244_0;
  wire [2:0] v_6245_0;
  wire [2:0] v_6246_0;
  wire [2:0] v_6247_0;
  reg [2:0] v_6248_0 = 3'h0;
  wire [0:0] v_6249_0;
  wire [0:0] v_6250_0;
  wire [0:0] v_6251_0;
  wire [2:0] v_6252_0;
  wire [2:0] v_6253_0;
  wire [2:0] v_6254_0;
  reg [2:0] v_6255_0 = 3'h0;
  wire [0:0] v_6256_0;
  wire [0:0] v_6257_0;
  wire [0:0] v_6258_0;
  wire [2:0] v_6259_0;
  wire [2:0] v_6260_0;
  wire [2:0] v_6261_0;
  reg [2:0] v_6262_0 = 3'h0;
  wire [0:0] v_6263_0;
  wire [0:0] v_6264_0;
  wire [0:0] v_6265_0;
  wire [2:0] v_6266_0;
  wire [2:0] v_6267_0;
  wire [2:0] v_6268_0;
  reg [2:0] v_6269_0 = 3'h0;
  wire [0:0] v_6270_0;
  wire [0:0] v_6271_0;
  wire [0:0] v_6272_0;
  wire [2:0] v_6273_0;
  wire [2:0] v_6274_0;
  wire [2:0] v_6275_0;
  reg [2:0] v_6276_0 = 3'h0;
  wire [0:0] v_6277_0;
  wire [0:0] v_6278_0;
  wire [0:0] v_6279_0;
  wire [2:0] v_6280_0;
  wire [2:0] v_6281_0;
  wire [2:0] v_6282_0;
  reg [2:0] v_6283_0 = 3'h0;
  wire [0:0] v_6284_0;
  wire [0:0] v_6285_0;
  wire [0:0] v_6286_0;
  wire [2:0] v_6287_0;
  wire [2:0] v_6288_0;
  wire [2:0] v_6289_0;
  reg [2:0] v_6290_0 = 3'h0;
  wire [0:0] v_6291_0;
  wire [0:0] v_6292_0;
  wire [0:0] v_6293_0;
  wire [2:0] v_6294_0;
  wire [2:0] v_6295_0;
  wire [2:0] v_6296_0;
  reg [2:0] v_6297_0 = 3'h0;
  wire [0:0] v_6298_0;
  wire [0:0] v_6299_0;
  wire [0:0] v_6300_0;
  wire [2:0] v_6301_0;
  wire [2:0] v_6302_0;
  wire [2:0] v_6303_0;
  reg [2:0] v_6304_0 = 3'h0;
  wire [0:0] v_6305_0;
  wire [0:0] v_6306_0;
  wire [0:0] v_6307_0;
  wire [2:0] v_6308_0;
  wire [2:0] v_6309_0;
  wire [2:0] v_6310_0;
  reg [2:0] v_6311_0 = 3'h0;
  wire [0:0] v_6312_0;
  wire [0:0] v_6313_0;
  wire [0:0] v_6314_0;
  wire [2:0] v_6315_0;
  wire [2:0] v_6316_0;
  wire [2:0] v_6317_0;
  reg [2:0] v_6318_0 = 3'h0;
  wire [0:0] v_6319_0;
  wire [0:0] v_6320_0;
  wire [0:0] v_6321_0;
  wire [2:0] v_6322_0;
  wire [2:0] v_6323_0;
  wire [2:0] v_6324_0;
  reg [2:0] v_6325_0 = 3'h0;
  wire [0:0] v_6326_0;
  wire [0:0] v_6327_0;
  wire [0:0] v_6328_0;
  wire [2:0] v_6329_0;
  wire [2:0] v_6330_0;
  wire [2:0] v_6331_0;
  reg [2:0] v_6332_0 = 3'h0;
  wire [0:0] v_6333_0;
  wire [0:0] v_6334_0;
  wire [0:0] v_6335_0;
  wire [2:0] v_6336_0;
  wire [2:0] v_6337_0;
  wire [2:0] v_6338_0;
  reg [2:0] v_6339_0 = 3'h0;
  wire [0:0] v_6340_0;
  wire [0:0] v_6341_0;
  wire [0:0] v_6342_0;
  wire [2:0] v_6343_0;
  wire [2:0] v_6344_0;
  wire [2:0] v_6345_0;
  reg [2:0] v_6346_0 = 3'h0;
  wire [0:0] v_6347_0;
  wire [0:0] v_6348_0;
  wire [0:0] v_6349_0;
  wire [2:0] v_6350_0;
  wire [2:0] v_6351_0;
  wire [2:0] v_6352_0;
  reg [2:0] v_6353_0 = 3'h0;
  wire [0:0] v_6354_0;
  wire [0:0] v_6355_0;
  wire [0:0] v_6356_0;
  wire [2:0] v_6357_0;
  wire [2:0] v_6358_0;
  wire [2:0] v_6359_0;
  reg [2:0] v_6360_0 = 3'h0;
  wire [0:0] v_6361_0;
  wire [0:0] v_6362_0;
  wire [0:0] v_6363_0;
  wire [2:0] v_6364_0;
  wire [2:0] v_6365_0;
  wire [2:0] v_6366_0;
  reg [2:0] v_6367_0 = 3'h0;
  wire [0:0] v_6368_0;
  wire [0:0] v_6369_0;
  wire [0:0] v_6370_0;
  wire [2:0] v_6371_0;
  wire [2:0] v_6372_0;
  wire [2:0] v_6373_0;
  reg [2:0] v_6374_0 = 3'h0;
  wire [0:0] v_6375_0;
  wire [0:0] v_6376_0;
  wire [0:0] v_6377_0;
  wire [2:0] v_6378_0;
  wire [2:0] v_6379_0;
  wire [2:0] v_6380_0;
  reg [2:0] v_6381_0 = 3'h0;
  wire [0:0] v_6382_0;
  wire [0:0] v_6383_0;
  wire [0:0] v_6384_0;
  wire [2:0] v_6385_0;
  wire [2:0] v_6386_0;
  wire [2:0] v_6387_0;
  reg [2:0] v_6388_0 = 3'h0;
  wire [0:0] v_6389_0;
  wire [0:0] v_6390_0;
  wire [0:0] v_6391_0;
  wire [2:0] v_6392_0;
  wire [2:0] v_6393_0;
  wire [2:0] v_6394_0;
  reg [2:0] v_6395_0 = 3'h0;
  wire [0:0] v_6396_0;
  wire [0:0] v_6397_0;
  wire [0:0] v_6398_0;
  wire [2:0] v_6399_0;
  wire [2:0] v_6400_0;
  wire [2:0] v_6401_0;
  reg [2:0] v_6402_0 = 3'h0;
  wire [0:0] v_6403_0;
  wire [0:0] v_6404_0;
  wire [0:0] v_6405_0;
  wire [2:0] v_6406_0;
  wire [2:0] v_6407_0;
  wire [2:0] v_6408_0;
  reg [2:0] v_6409_0 = 3'h0;
  wire [0:0] v_6410_0;
  wire [0:0] v_6411_0;
  wire [0:0] v_6412_0;
  wire [2:0] v_6413_0;
  wire [2:0] v_6414_0;
  wire [2:0] v_6415_0;
  reg [2:0] v_6416_0 = 3'h0;
  wire [0:0] v_6417_0;
  wire [0:0] v_6418_0;
  wire [0:0] v_6419_0;
  wire [2:0] v_6420_0;
  wire [2:0] v_6421_0;
  wire [2:0] v_6422_0;
  reg [2:0] v_6423_0 = 3'h0;
  wire [0:0] v_6424_0;
  wire [0:0] v_6425_0;
  wire [0:0] v_6426_0;
  wire [2:0] v_6427_0;
  wire [2:0] v_6428_0;
  wire [2:0] v_6429_0;
  reg [2:0] v_6430_0 = 3'h0;
  wire [0:0] v_6431_0;
  wire [0:0] v_6432_0;
  wire [0:0] v_6433_0;
  wire [2:0] v_6434_0;
  wire [2:0] v_6435_0;
  wire [2:0] v_6436_0;
  reg [2:0] v_6437_0 = 3'h0;
  wire [0:0] v_6438_0;
  wire [0:0] v_6439_0;
  wire [0:0] v_6440_0;
  wire [2:0] v_6441_0;
  wire [2:0] v_6442_0;
  wire [2:0] v_6443_0;
  reg [2:0] v_6444_0 = 3'h0;
  wire [0:0] v_6445_0;
  wire [0:0] v_6446_0;
  wire [0:0] v_6447_0;
  wire [2:0] v_6448_0;
  wire [2:0] v_6449_0;
  wire [2:0] v_6450_0;
  reg [2:0] v_6451_0 = 3'h0;
  wire [0:0] v_6452_0;
  wire [0:0] v_6453_0;
  wire [0:0] v_6454_0;
  wire [2:0] v_6455_0;
  wire [2:0] v_6456_0;
  wire [2:0] v_6457_0;
  reg [2:0] v_6458_0 = 3'h0;
  wire [0:0] v_6459_0;
  wire [0:0] v_6460_0;
  wire [0:0] v_6461_0;
  wire [2:0] v_6462_0;
  wire [2:0] v_6463_0;
  wire [2:0] v_6464_0;
  reg [2:0] v_6465_0 = 3'h0;
  wire [0:0] v_6466_0;
  wire [0:0] v_6467_0;
  wire [0:0] v_6468_0;
  wire [2:0] v_6469_0;
  wire [2:0] v_6470_0;
  wire [2:0] v_6471_0;
  reg [2:0] v_6472_0 = 3'h0;
  wire [0:0] v_6473_0;
  wire [0:0] v_6474_0;
  wire [0:0] v_6475_0;
  wire [2:0] v_6476_0;
  wire [2:0] v_6477_0;
  wire [2:0] v_6478_0;
  reg [2:0] v_6479_0 = 3'h0;
  wire [0:0] v_6480_0;
  wire [0:0] v_6481_0;
  wire [0:0] v_6482_0;
  wire [2:0] v_6483_0;
  wire [2:0] v_6484_0;
  wire [2:0] v_6485_0;
  reg [2:0] v_6486_0 = 3'h0;
  wire [0:0] v_6487_0;
  wire [0:0] v_6488_0;
  wire [0:0] v_6489_0;
  wire [2:0] v_6490_0;
  wire [2:0] v_6491_0;
  wire [2:0] v_6492_0;
  reg [2:0] v_6493_0 = 3'h0;
  wire [0:0] v_6494_0;
  wire [0:0] v_6495_0;
  wire [0:0] v_6496_0;
  wire [2:0] v_6497_0;
  wire [2:0] v_6498_0;
  wire [2:0] v_6499_0;
  reg [2:0] v_6500_0 = 3'h0;
  wire [0:0] v_6501_0;
  wire [0:0] v_6502_0;
  wire [0:0] v_6503_0;
  wire [2:0] v_6504_0;
  wire [2:0] v_6505_0;
  wire [2:0] v_6506_0;
  reg [2:0] v_6507_0 = 3'h0;
  wire [0:0] v_6508_0;
  wire [0:0] v_6509_0;
  wire [0:0] v_6510_0;
  wire [2:0] v_6511_0;
  wire [2:0] v_6512_0;
  wire [2:0] v_6513_0;
  reg [2:0] v_6514_0 = 3'h0;
  wire [0:0] v_6515_0;
  wire [0:0] v_6516_0;
  wire [0:0] v_6517_0;
  wire [2:0] v_6518_0;
  wire [2:0] v_6519_0;
  wire [2:0] v_6520_0;
  reg [2:0] v_6521_0 = 3'h0;
  wire [0:0] v_6522_0;
  wire [0:0] v_6523_0;
  wire [0:0] v_6524_0;
  wire [2:0] v_6525_0;
  wire [2:0] v_6526_0;
  wire [2:0] v_6527_0;
  reg [2:0] v_6528_0 = 3'h0;
  wire [0:0] v_6529_0;
  wire [0:0] v_6530_0;
  wire [0:0] v_6531_0;
  wire [2:0] v_6532_0;
  wire [2:0] v_6533_0;
  wire [2:0] v_6534_0;
  reg [2:0] v_6535_0 = 3'h0;
  wire [0:0] v_6536_0;
  wire [0:0] v_6537_0;
  wire [0:0] v_6538_0;
  wire [2:0] v_6539_0;
  wire [2:0] v_6540_0;
  wire [2:0] v_6541_0;
  reg [2:0] v_6542_0 = 3'h0;
  wire [0:0] v_6543_0;
  wire [0:0] v_6544_0;
  wire [0:0] v_6545_0;
  wire [2:0] v_6546_0;
  wire [2:0] v_6547_0;
  wire [2:0] v_6548_0;
  reg [2:0] v_6549_0 = 3'h0;
  wire [0:0] v_6550_0;
  wire [0:0] v_6551_0;
  wire [0:0] v_6552_0;
  wire [2:0] v_6553_0;
  wire [2:0] v_6554_0;
  wire [2:0] v_6555_0;
  reg [2:0] v_6556_0 = 3'h0;
  wire [0:0] v_6557_0;
  wire [0:0] v_6558_0;
  wire [0:0] v_6559_0;
  wire [2:0] v_6560_0;
  wire [2:0] v_6561_0;
  wire [2:0] v_6562_0;
  reg [2:0] v_6563_0 = 3'h0;
  wire [0:0] v_6564_0;
  wire [0:0] v_6565_0;
  wire [0:0] v_6566_0;
  wire [2:0] v_6567_0;
  wire [2:0] v_6568_0;
  wire [2:0] v_6569_0;
  reg [2:0] v_6570_0 = 3'h0;
  wire [0:0] v_6571_0;
  wire [0:0] v_6572_0;
  wire [0:0] v_6573_0;
  wire [2:0] v_6574_0;
  wire [2:0] v_6575_0;
  wire [2:0] v_6576_0;
  reg [2:0] v_6577_0 = 3'h0;
  wire [0:0] v_6578_0;
  wire [0:0] v_6579_0;
  wire [0:0] v_6580_0;
  wire [2:0] v_6581_0;
  wire [2:0] v_6582_0;
  wire [2:0] v_6583_0;
  reg [2:0] v_6584_0 = 3'h0;
  wire [0:0] v_6585_0;
  wire [0:0] v_6586_0;
  wire [0:0] v_6587_0;
  wire [2:0] v_6588_0;
  wire [2:0] v_6589_0;
  wire [2:0] v_6590_0;
  reg [2:0] v_6591_0 = 3'h0;
  wire [0:0] v_6592_0;
  wire [0:0] v_6593_0;
  wire [0:0] v_6594_0;
  wire [2:0] v_6595_0;
  wire [2:0] v_6596_0;
  wire [2:0] v_6597_0;
  reg [2:0] v_6598_0 = 3'h0;
  wire [0:0] v_6599_0;
  wire [0:0] v_6600_0;
  wire [0:0] v_6601_0;
  wire [2:0] v_6602_0;
  wire [2:0] v_6603_0;
  wire [2:0] v_6604_0;
  reg [2:0] v_6605_0 = 3'h0;
  wire [0:0] v_6606_0;
  wire [0:0] v_6607_0;
  wire [0:0] v_6608_0;
  wire [2:0] v_6609_0;
  wire [2:0] v_6610_0;
  wire [2:0] v_6611_0;
  reg [2:0] v_6612_0 = 3'h0;
  wire [0:0] v_6613_0;
  wire [0:0] v_6614_0;
  wire [0:0] v_6615_0;
  wire [2:0] v_6616_0;
  wire [2:0] v_6617_0;
  wire [2:0] v_6618_0;
  reg [2:0] v_6619_0 = 3'h0;
  wire [0:0] v_6620_0;
  wire [0:0] v_6621_0;
  wire [0:0] v_6622_0;
  wire [2:0] v_6623_0;
  wire [2:0] v_6624_0;
  wire [2:0] v_6625_0;
  reg [2:0] v_6626_0 = 3'h0;
  wire [0:0] v_6627_0;
  wire [0:0] v_6628_0;
  wire [0:0] v_6629_0;
  wire [2:0] v_6630_0;
  wire [2:0] v_6631_0;
  wire [2:0] v_6632_0;
  reg [2:0] v_6633_0 = 3'h0;
  wire [0:0] v_6634_0;
  wire [0:0] v_6635_0;
  wire [0:0] v_6636_0;
  wire [2:0] v_6637_0;
  wire [2:0] v_6638_0;
  wire [2:0] v_6639_0;
  reg [2:0] v_6640_0 = 3'h0;
  wire [0:0] v_6641_0;
  wire [0:0] v_6642_0;
  wire [0:0] v_6643_0;
  wire [2:0] v_6644_0;
  wire [2:0] v_6645_0;
  wire [2:0] v_6646_0;
  reg [2:0] v_6647_0 = 3'h0;
  wire [0:0] v_6648_0;
  wire [0:0] v_6649_0;
  wire [0:0] v_6650_0;
  wire [2:0] v_6651_0;
  wire [2:0] v_6652_0;
  wire [2:0] v_6653_0;
  reg [2:0] v_6654_0 = 3'h0;
  wire [0:0] v_6655_0;
  wire [0:0] v_6656_0;
  wire [0:0] v_6657_0;
  wire [2:0] v_6658_0;
  wire [2:0] v_6659_0;
  wire [2:0] v_6660_0;
  reg [2:0] v_6661_0 = 3'h0;
  wire [0:0] v_6662_0;
  wire [0:0] v_6663_0;
  wire [0:0] v_6664_0;
  wire [2:0] v_6665_0;
  wire [2:0] v_6666_0;
  wire [2:0] v_6667_0;
  reg [2:0] v_6668_0 = 3'h0;
  wire [0:0] v_6669_0;
  wire [0:0] v_6670_0;
  wire [0:0] v_6671_0;
  wire [2:0] v_6672_0;
  wire [2:0] v_6673_0;
  wire [2:0] v_6674_0;
  reg [2:0] v_6675_0 = 3'h0;
  wire [0:0] v_6676_0;
  wire [0:0] v_6677_0;
  wire [0:0] v_6678_0;
  wire [2:0] v_6679_0;
  wire [2:0] v_6680_0;
  wire [2:0] v_6681_0;
  reg [2:0] v_6682_0 = 3'h0;
  wire [0:0] v_6683_0;
  wire [0:0] v_6684_0;
  wire [0:0] v_6685_0;
  wire [2:0] v_6686_0;
  wire [2:0] v_6687_0;
  wire [2:0] v_6688_0;
  reg [2:0] v_6689_0 = 3'h0;
  wire [0:0] v_6690_0;
  wire [0:0] v_6691_0;
  wire [0:0] v_6692_0;
  wire [2:0] v_6693_0;
  wire [2:0] v_6694_0;
  wire [2:0] v_6695_0;
  reg [2:0] v_6696_0 = 3'h0;
  wire [0:0] v_6697_0;
  wire [0:0] v_6698_0;
  wire [0:0] v_6699_0;
  wire [2:0] v_6700_0;
  wire [2:0] v_6701_0;
  wire [2:0] v_6702_0;
  reg [2:0] v_6703_0 = 3'h0;
  wire [0:0] v_6704_0;
  wire [0:0] v_6705_0;
  wire [0:0] v_6706_0;
  wire [2:0] v_6707_0;
  wire [2:0] v_6708_0;
  wire [2:0] v_6709_0;
  reg [2:0] v_6710_0 = 3'h0;
  wire [0:0] v_6711_0;
  wire [0:0] v_6712_0;
  wire [0:0] v_6713_0;
  wire [2:0] v_6714_0;
  wire [2:0] v_6715_0;
  wire [2:0] v_6716_0;
  reg [2:0] v_6717_0 = 3'h0;
  wire [0:0] v_6718_0;
  wire [0:0] v_6719_0;
  wire [0:0] v_6720_0;
  wire [2:0] v_6721_0;
  wire [2:0] v_6722_0;
  wire [2:0] v_6723_0;
  reg [2:0] v_6724_0 = 3'h0;
  wire [0:0] v_6725_0;
  wire [0:0] v_6726_0;
  wire [0:0] v_6727_0;
  wire [2:0] v_6728_0;
  wire [2:0] v_6729_0;
  wire [2:0] v_6730_0;
  reg [2:0] v_6731_0 = 3'h0;
  wire [0:0] v_6732_0;
  wire [0:0] v_6733_0;
  wire [0:0] v_6734_0;
  wire [2:0] v_6735_0;
  wire [2:0] v_6736_0;
  wire [2:0] v_6737_0;
  reg [2:0] v_6738_0 = 3'h0;
  wire [0:0] v_6739_0;
  wire [0:0] v_6740_0;
  wire [0:0] v_6741_0;
  wire [2:0] v_6742_0;
  wire [2:0] v_6743_0;
  wire [2:0] v_6744_0;
  reg [2:0] v_6745_0 = 3'h0;
  wire [0:0] v_6746_0;
  wire [0:0] v_6747_0;
  wire [0:0] v_6748_0;
  wire [2:0] v_6749_0;
  wire [2:0] v_6750_0;
  wire [2:0] v_6751_0;
  reg [2:0] v_6752_0 = 3'h0;
  wire [0:0] v_6753_0;
  wire [0:0] v_6754_0;
  wire [0:0] v_6755_0;
  wire [2:0] v_6756_0;
  wire [2:0] v_6757_0;
  wire [2:0] v_6758_0;
  reg [2:0] v_6759_0 = 3'h0;
  wire [0:0] v_6760_0;
  wire [0:0] v_6761_0;
  wire [0:0] v_6762_0;
  wire [2:0] v_6763_0;
  wire [2:0] v_6764_0;
  wire [2:0] v_6765_0;
  reg [2:0] v_6766_0 = 3'h0;
  wire [0:0] v_6767_0;
  wire [0:0] v_6768_0;
  wire [0:0] v_6769_0;
  wire [2:0] v_6770_0;
  wire [2:0] v_6771_0;
  wire [2:0] v_6772_0;
  reg [2:0] v_6773_0 = 3'h0;
  wire [0:0] v_6774_0;
  wire [0:0] v_6775_0;
  wire [0:0] v_6776_0;
  wire [2:0] v_6777_0;
  wire [2:0] v_6778_0;
  wire [2:0] v_6779_0;
  reg [2:0] v_6780_0 = 3'h0;
  wire [0:0] v_6781_0;
  wire [0:0] v_6782_0;
  wire [0:0] v_6783_0;
  wire [2:0] v_6784_0;
  wire [2:0] v_6785_0;
  wire [2:0] v_6786_0;
  reg [2:0] v_6787_0 = 3'h0;
  wire [0:0] v_6788_0;
  wire [0:0] v_6789_0;
  wire [0:0] v_6790_0;
  wire [2:0] v_6791_0;
  wire [2:0] v_6792_0;
  wire [2:0] v_6793_0;
  reg [2:0] v_6794_0 = 3'h0;
  wire [0:0] v_6795_0;
  wire [0:0] v_6796_0;
  wire [0:0] v_6797_0;
  wire [2:0] v_6798_0;
  wire [2:0] v_6799_0;
  wire [2:0] v_6800_0;
  reg [2:0] v_6801_0 = 3'h0;
  wire [0:0] v_6802_0;
  wire [0:0] v_6803_0;
  wire [0:0] v_6804_0;
  wire [2:0] v_6805_0;
  wire [2:0] v_6806_0;
  wire [2:0] v_6807_0;
  reg [2:0] v_6808_0 = 3'h0;
  wire [0:0] v_6809_0;
  wire [0:0] v_6810_0;
  wire [0:0] v_6811_0;
  wire [2:0] v_6812_0;
  wire [2:0] v_6813_0;
  wire [2:0] v_6814_0;
  reg [2:0] v_6815_0 = 3'h0;
  wire [0:0] v_6816_0;
  wire [0:0] v_6817_0;
  wire [0:0] v_6818_0;
  wire [2:0] v_6819_0;
  wire [2:0] v_6820_0;
  wire [2:0] v_6821_0;
  reg [2:0] v_6822_0 = 3'h0;
  wire [0:0] v_6823_0;
  wire [0:0] v_6824_0;
  wire [0:0] v_6825_0;
  wire [2:0] v_6826_0;
  wire [2:0] v_6827_0;
  wire [2:0] v_6828_0;
  reg [2:0] v_6829_0 = 3'h0;
  wire [0:0] v_6830_0;
  wire [0:0] v_6831_0;
  wire [0:0] v_6832_0;
  wire [2:0] v_6833_0;
  wire [2:0] v_6834_0;
  wire [2:0] v_6835_0;
  reg [2:0] v_6836_0 = 3'h0;
  wire [0:0] v_6837_0;
  wire [0:0] v_6838_0;
  wire [0:0] v_6839_0;
  wire [2:0] v_6840_0;
  wire [2:0] v_6841_0;
  wire [2:0] v_6842_0;
  reg [2:0] v_6843_0 = 3'h0;
  wire [0:0] v_6844_0;
  wire [0:0] v_6845_0;
  wire [0:0] v_6846_0;
  wire [2:0] v_6847_0;
  wire [2:0] v_6848_0;
  wire [2:0] v_6849_0;
  reg [2:0] v_6850_0 = 3'h0;
  wire [0:0] v_6851_0;
  wire [0:0] v_6852_0;
  wire [0:0] v_6853_0;
  wire [2:0] v_6854_0;
  wire [2:0] v_6855_0;
  wire [2:0] v_6856_0;
  reg [2:0] v_6857_0 = 3'h0;
  wire [0:0] v_6858_0;
  wire [0:0] v_6859_0;
  wire [0:0] v_6860_0;
  wire [2:0] v_6861_0;
  wire [2:0] v_6862_0;
  wire [2:0] v_6863_0;
  reg [2:0] v_6864_0 = 3'h0;
  wire [0:0] v_6865_0;
  wire [0:0] v_6866_0;
  wire [0:0] v_6867_0;
  wire [2:0] v_6868_0;
  wire [2:0] v_6869_0;
  wire [2:0] v_6870_0;
  reg [2:0] v_6871_0 = 3'h0;
  wire [0:0] v_6872_0;
  wire [0:0] v_6873_0;
  wire [0:0] v_6874_0;
  wire [2:0] v_6875_0;
  wire [2:0] v_6876_0;
  wire [2:0] v_6877_0;
  reg [2:0] v_6878_0 = 3'h0;
  wire [0:0] v_6879_0;
  wire [0:0] v_6880_0;
  wire [0:0] v_6881_0;
  wire [2:0] v_6882_0;
  wire [2:0] v_6883_0;
  wire [2:0] v_6884_0;
  reg [2:0] v_6885_0 = 3'h0;
  wire [0:0] v_6886_0;
  wire [0:0] v_6887_0;
  wire [0:0] v_6888_0;
  wire [2:0] v_6889_0;
  wire [2:0] v_6890_0;
  wire [2:0] v_6891_0;
  reg [2:0] v_6892_0 = 3'h0;
  wire [0:0] v_6893_0;
  wire [0:0] v_6894_0;
  wire [0:0] v_6895_0;
  wire [2:0] v_6896_0;
  wire [2:0] v_6897_0;
  wire [2:0] v_6898_0;
  reg [2:0] v_6899_0 = 3'h0;
  wire [0:0] v_6900_0;
  wire [0:0] v_6901_0;
  wire [0:0] v_6902_0;
  wire [2:0] v_6903_0;
  wire [2:0] v_6904_0;
  wire [2:0] v_6905_0;
  reg [2:0] v_6906_0 = 3'h0;
  wire [0:0] v_6907_0;
  wire [0:0] v_6908_0;
  wire [0:0] v_6909_0;
  wire [2:0] v_6910_0;
  wire [2:0] v_6911_0;
  wire [2:0] v_6912_0;
  reg [2:0] v_6913_0 = 3'h0;
  wire [0:0] v_6914_0;
  wire [0:0] v_6915_0;
  wire [0:0] v_6916_0;
  wire [2:0] v_6917_0;
  wire [2:0] v_6918_0;
  wire [2:0] v_6919_0;
  reg [2:0] v_6920_0 = 3'h0;
  wire [0:0] v_6921_0;
  wire [0:0] v_6922_0;
  wire [0:0] v_6923_0;
  wire [2:0] v_6924_0;
  wire [2:0] v_6925_0;
  wire [2:0] v_6926_0;
  reg [2:0] v_6927_0 = 3'h0;
  wire [0:0] v_6928_0;
  wire [0:0] v_6929_0;
  wire [0:0] v_6930_0;
  wire [2:0] v_6931_0;
  wire [2:0] v_6932_0;
  wire [2:0] v_6933_0;
  reg [2:0] v_6934_0 = 3'h0;
  wire [0:0] v_6935_0;
  wire [0:0] v_6936_0;
  wire [0:0] v_6937_0;
  wire [2:0] v_6938_0;
  wire [2:0] v_6939_0;
  wire [2:0] v_6940_0;
  reg [2:0] v_6941_0 = 3'h0;
  wire [0:0] v_6942_0;
  wire [0:0] v_6943_0;
  wire [0:0] v_6944_0;
  wire [2:0] v_6945_0;
  wire [2:0] v_6946_0;
  wire [2:0] v_6947_0;
  reg [2:0] v_6948_0 = 3'h0;
  wire [0:0] v_6949_0;
  wire [0:0] v_6950_0;
  wire [0:0] v_6951_0;
  wire [2:0] v_6952_0;
  wire [2:0] v_6953_0;
  wire [2:0] v_6954_0;
  reg [2:0] v_6955_0 = 3'h0;
  wire [0:0] v_6956_0;
  wire [0:0] v_6957_0;
  wire [0:0] v_6958_0;
  wire [2:0] v_6959_0;
  wire [2:0] v_6960_0;
  wire [2:0] v_6961_0;
  reg [2:0] v_6962_0 = 3'h0;
  wire [0:0] v_6963_0;
  wire [0:0] v_6964_0;
  wire [0:0] v_6965_0;
  wire [2:0] v_6966_0;
  wire [2:0] v_6967_0;
  wire [2:0] v_6968_0;
  reg [2:0] v_6969_0 = 3'h0;
  wire [0:0] v_6970_0;
  wire [0:0] v_6971_0;
  wire [0:0] v_6972_0;
  wire [2:0] v_6973_0;
  wire [2:0] v_6974_0;
  wire [2:0] v_6975_0;
  reg [2:0] v_6976_0 = 3'h0;
  wire [0:0] v_6977_0;
  wire [0:0] v_6978_0;
  wire [0:0] v_6979_0;
  wire [2:0] v_6980_0;
  wire [2:0] v_6981_0;
  wire [2:0] v_6982_0;
  reg [2:0] v_6983_0 = 3'h0;
  wire [0:0] v_6984_0;
  wire [0:0] v_6985_0;
  wire [0:0] v_6986_0;
  wire [2:0] v_6987_0;
  wire [2:0] v_6988_0;
  wire [2:0] v_6989_0;
  reg [2:0] v_6990_0 = 3'h0;
  wire [0:0] v_6991_0;
  wire [0:0] v_6992_0;
  wire [0:0] v_6993_0;
  wire [2:0] v_6994_0;
  wire [2:0] v_6995_0;
  wire [2:0] v_6996_0;
  reg [2:0] v_6997_0 = 3'h0;
  wire [0:0] v_6998_0;
  wire [0:0] v_6999_0;
  wire [0:0] v_7000_0;
  wire [2:0] v_7001_0;
  wire [2:0] v_7002_0;
  wire [2:0] v_7003_0;
  reg [2:0] v_7004_0 = 3'h0;
  wire [0:0] v_7005_0;
  wire [0:0] v_7006_0;
  wire [0:0] v_7007_0;
  wire [2:0] v_7008_0;
  wire [2:0] v_7009_0;
  wire [2:0] v_7010_0;
  reg [2:0] v_7011_0 = 3'h0;
  wire [0:0] v_7012_0;
  wire [0:0] v_7013_0;
  wire [0:0] v_7014_0;
  wire [2:0] v_7015_0;
  wire [2:0] v_7016_0;
  wire [2:0] v_7017_0;
  reg [2:0] v_7018_0 = 3'h0;
  wire [0:0] v_7019_0;
  wire [0:0] v_7020_0;
  wire [0:0] v_7021_0;
  wire [2:0] v_7022_0;
  wire [2:0] v_7023_0;
  wire [2:0] v_7024_0;
  reg [2:0] v_7025_0 = 3'h0;
  wire [0:0] v_7026_0;
  wire [0:0] v_7027_0;
  wire [0:0] v_7028_0;
  wire [2:0] v_7029_0;
  wire [2:0] v_7030_0;
  wire [2:0] v_7031_0;
  reg [2:0] v_7032_0 = 3'h0;
  wire [0:0] v_7033_0;
  wire [0:0] v_7034_0;
  wire [0:0] v_7035_0;
  wire [2:0] v_7036_0;
  wire [2:0] v_7037_0;
  wire [2:0] v_7038_0;
  reg [2:0] v_7039_0 = 3'h0;
  wire [0:0] v_7040_0;
  wire [0:0] v_7041_0;
  wire [0:0] v_7042_0;
  wire [2:0] v_7043_0;
  wire [2:0] v_7044_0;
  wire [2:0] v_7045_0;
  reg [2:0] v_7046_0 = 3'h0;
  wire [0:0] v_7047_0;
  wire [0:0] v_7048_0;
  wire [0:0] v_7049_0;
  wire [2:0] v_7050_0;
  wire [2:0] v_7051_0;
  wire [2:0] v_7052_0;
  reg [2:0] v_7053_0 = 3'h0;
  wire [0:0] v_7054_0;
  wire [0:0] v_7055_0;
  wire [0:0] v_7056_0;
  wire [2:0] v_7057_0;
  wire [2:0] v_7058_0;
  wire [2:0] v_7059_0;
  reg [2:0] v_7060_0 = 3'h0;
  wire [0:0] v_7061_0;
  wire [0:0] v_7062_0;
  wire [0:0] v_7063_0;
  wire [2:0] v_7064_0;
  wire [2:0] v_7065_0;
  wire [2:0] v_7066_0;
  reg [2:0] v_7067_0 = 3'h0;
  wire [0:0] v_7068_0;
  wire [0:0] v_7069_0;
  wire [0:0] v_7070_0;
  wire [2:0] v_7071_0;
  wire [2:0] v_7072_0;
  wire [2:0] v_7073_0;
  reg [2:0] v_7074_0 = 3'h0;
  wire [0:0] v_7075_0;
  wire [0:0] v_7076_0;
  wire [0:0] v_7077_0;
  wire [2:0] v_7078_0;
  wire [2:0] v_7079_0;
  wire [2:0] v_7080_0;
  reg [2:0] v_7081_0 = 3'h0;
  wire [0:0] v_7082_0;
  wire [0:0] v_7083_0;
  wire [0:0] v_7084_0;
  wire [2:0] v_7085_0;
  wire [2:0] v_7086_0;
  wire [2:0] v_7087_0;
  reg [2:0] v_7088_0 = 3'h0;
  wire [0:0] v_7089_0;
  wire [0:0] v_7090_0;
  wire [0:0] v_7091_0;
  wire [2:0] v_7092_0;
  wire [2:0] v_7093_0;
  wire [2:0] v_7094_0;
  reg [2:0] v_7095_0 = 3'h0;
  wire [0:0] v_7096_0;
  wire [0:0] v_7097_0;
  wire [0:0] v_7098_0;
  wire [2:0] v_7099_0;
  wire [2:0] v_7100_0;
  wire [2:0] v_7101_0;
  reg [2:0] v_7102_0 = 3'h0;
  wire [0:0] v_7103_0;
  wire [0:0] v_7104_0;
  wire [0:0] v_7105_0;
  wire [2:0] v_7106_0;
  wire [2:0] v_7107_0;
  wire [2:0] v_7108_0;
  reg [2:0] v_7109_0 = 3'h0;
  wire [0:0] v_7110_0;
  wire [0:0] v_7111_0;
  wire [0:0] v_7112_0;
  wire [2:0] v_7113_0;
  wire [2:0] v_7114_0;
  wire [2:0] v_7115_0;
  reg [2:0] v_7116_0 = 3'h0;
  wire [0:0] v_7117_0;
  wire [0:0] v_7118_0;
  wire [0:0] v_7119_0;
  wire [2:0] v_7120_0;
  wire [2:0] v_7121_0;
  wire [2:0] v_7122_0;
  reg [2:0] v_7123_0 = 3'h0;
  wire [0:0] v_7124_0;
  wire [0:0] v_7125_0;
  wire [0:0] v_7126_0;
  wire [2:0] v_7127_0;
  wire [2:0] v_7128_0;
  wire [2:0] v_7129_0;
  reg [2:0] v_7130_0 = 3'h0;
  wire [0:0] v_7131_0;
  wire [0:0] v_7132_0;
  wire [0:0] v_7133_0;
  wire [2:0] v_7134_0;
  wire [2:0] v_7135_0;
  wire [2:0] v_7136_0;
  reg [2:0] v_7137_0 = 3'h0;
  wire [0:0] v_7138_0;
  wire [0:0] v_7139_0;
  wire [0:0] v_7140_0;
  wire [2:0] v_7141_0;
  wire [2:0] v_7142_0;
  wire [2:0] v_7143_0;
  reg [2:0] v_7144_0 = 3'h0;
  wire [0:0] v_7145_0;
  wire [0:0] v_7146_0;
  wire [0:0] v_7147_0;
  wire [2:0] v_7148_0;
  wire [2:0] v_7149_0;
  wire [2:0] v_7150_0;
  reg [2:0] v_7151_0 = 3'h0;
  wire [0:0] v_7152_0;
  wire [0:0] v_7153_0;
  wire [0:0] v_7154_0;
  wire [2:0] v_7155_0;
  wire [2:0] v_7156_0;
  wire [2:0] v_7157_0;
  reg [2:0] v_7158_0 = 3'h0;
  wire [0:0] v_7159_0;
  wire [0:0] v_7160_0;
  wire [0:0] v_7161_0;
  wire [2:0] v_7162_0;
  wire [2:0] v_7163_0;
  wire [2:0] v_7164_0;
  reg [2:0] v_7165_0 = 3'h0;
  wire [0:0] v_7166_0;
  wire [0:0] v_7167_0;
  wire [0:0] v_7168_0;
  wire [2:0] v_7169_0;
  wire [2:0] v_7170_0;
  wire [2:0] v_7171_0;
  reg [2:0] v_7172_0 = 3'h0;
  wire [0:0] v_7173_0;
  wire [0:0] v_7174_0;
  wire [0:0] v_7175_0;
  wire [2:0] v_7176_0;
  wire [2:0] v_7177_0;
  wire [2:0] v_7178_0;
  reg [2:0] v_7179_0 = 3'h0;
  wire [0:0] v_7180_0;
  wire [0:0] v_7181_0;
  wire [0:0] v_7182_0;
  wire [2:0] v_7183_0;
  wire [2:0] v_7184_0;
  wire [2:0] v_7185_0;
  reg [2:0] v_7186_0 = 3'h0;
  wire [0:0] v_7187_0;
  wire [0:0] v_7188_0;
  wire [0:0] v_7189_0;
  wire [2:0] v_7190_0;
  wire [2:0] v_7191_0;
  wire [2:0] v_7192_0;
  reg [2:0] v_7193_0 = 3'h0;
  wire [0:0] v_7194_0;
  wire [0:0] v_7195_0;
  wire [0:0] v_7196_0;
  wire [2:0] v_7197_0;
  wire [2:0] v_7198_0;
  wire [2:0] v_7199_0;
  reg [2:0] v_7200_0 = 3'h0;
  wire [0:0] v_7201_0;
  wire [0:0] v_7202_0;
  wire [0:0] v_7203_0;
  wire [2:0] v_7204_0;
  wire [2:0] v_7205_0;
  wire [2:0] v_7206_0;
  reg [2:0] v_7207_0 = 3'h0;
  wire [0:0] v_7208_0;
  wire [0:0] v_7209_0;
  wire [0:0] v_7210_0;
  wire [2:0] v_7211_0;
  wire [2:0] v_7212_0;
  wire [2:0] v_7213_0;
  reg [2:0] v_7214_0 = 3'h0;
  wire [0:0] v_7215_0;
  wire [0:0] v_7216_0;
  wire [0:0] v_7217_0;
  wire [2:0] v_7218_0;
  wire [2:0] v_7219_0;
  wire [2:0] v_7220_0;
  reg [2:0] v_7221_0 = 3'h0;
  wire [0:0] v_7222_0;
  wire [0:0] v_7223_0;
  wire [0:0] v_7224_0;
  wire [2:0] v_7225_0;
  wire [2:0] v_7226_0;
  wire [2:0] v_7227_0;
  reg [2:0] v_7228_0 = 3'h0;
  wire [0:0] v_7229_0;
  wire [0:0] v_7230_0;
  wire [0:0] v_7231_0;
  wire [2:0] v_7232_0;
  wire [2:0] v_7233_0;
  wire [2:0] v_7234_0;
  reg [2:0] v_7235_0 = 3'h0;
  wire [0:0] v_7236_0;
  wire [0:0] v_7237_0;
  wire [0:0] v_7238_0;
  wire [2:0] v_7239_0;
  wire [2:0] v_7240_0;
  wire [2:0] v_7241_0;
  reg [2:0] v_7242_0 = 3'h0;
  wire [0:0] v_7243_0;
  wire [0:0] v_7244_0;
  wire [0:0] v_7245_0;
  wire [2:0] v_7246_0;
  wire [2:0] v_7247_0;
  wire [2:0] v_7248_0;
  reg [2:0] v_7249_0 = 3'h0;
  wire [0:0] v_7250_0;
  wire [0:0] v_7251_0;
  wire [0:0] v_7252_0;
  wire [2:0] v_7253_0;
  wire [2:0] v_7254_0;
  wire [2:0] v_7255_0;
  reg [2:0] v_7256_0 = 3'h0;
  wire [0:0] v_7257_0;
  wire [0:0] v_7258_0;
  wire [0:0] v_7259_0;
  wire [2:0] v_7260_0;
  wire [2:0] v_7261_0;
  wire [2:0] v_7262_0;
  reg [2:0] v_7263_0 = 3'h0;
  wire [0:0] v_7264_0;
  wire [0:0] v_7265_0;
  wire [0:0] v_7266_0;
  wire [2:0] v_7267_0;
  wire [2:0] v_7268_0;
  wire [2:0] v_7269_0;
  reg [2:0] v_7270_0 = 3'h0;
  wire [0:0] v_7271_0;
  wire [0:0] v_7272_0;
  wire [0:0] v_7273_0;
  wire [2:0] v_7274_0;
  wire [2:0] v_7275_0;
  wire [2:0] v_7276_0;
  reg [2:0] v_7277_0 = 3'h0;
  wire [0:0] v_7278_0;
  wire [0:0] v_7279_0;
  wire [0:0] v_7280_0;
  wire [2:0] v_7281_0;
  wire [2:0] v_7282_0;
  wire [2:0] v_7283_0;
  reg [2:0] v_7284_0 = 3'h0;
  wire [0:0] v_7285_0;
  wire [0:0] v_7286_0;
  wire [0:0] v_7287_0;
  wire [2:0] v_7288_0;
  wire [2:0] v_7289_0;
  wire [2:0] v_7290_0;
  reg [2:0] v_7291_0 = 3'h0;
  wire [0:0] v_7292_0;
  wire [0:0] v_7293_0;
  wire [0:0] v_7294_0;
  wire [2:0] v_7295_0;
  wire [2:0] v_7296_0;
  wire [2:0] v_7297_0;
  reg [2:0] v_7298_0 = 3'h0;
  wire [0:0] v_7299_0;
  wire [0:0] v_7300_0;
  wire [0:0] v_7301_0;
  wire [2:0] v_7302_0;
  wire [2:0] v_7303_0;
  wire [2:0] v_7304_0;
  reg [2:0] v_7305_0 = 3'h0;
  wire [0:0] v_7306_0;
  wire [0:0] v_7307_0;
  wire [0:0] v_7308_0;
  wire [2:0] v_7309_0;
  wire [2:0] v_7310_0;
  wire [2:0] v_7311_0;
  reg [2:0] v_7312_0 = 3'h0;
  wire [0:0] v_7313_0;
  wire [0:0] v_7314_0;
  wire [0:0] v_7315_0;
  wire [2:0] v_7316_0;
  wire [2:0] v_7317_0;
  wire [2:0] v_7318_0;
  reg [2:0] v_7319_0 = 3'h0;
  wire [0:0] v_7320_0;
  wire [0:0] v_7321_0;
  wire [0:0] v_7322_0;
  wire [2:0] v_7323_0;
  wire [2:0] v_7324_0;
  wire [2:0] v_7325_0;
  reg [2:0] v_7326_0 = 3'h0;
  wire [0:0] v_7327_0;
  wire [0:0] v_7328_0;
  wire [0:0] v_7329_0;
  wire [2:0] v_7330_0;
  wire [2:0] v_7331_0;
  wire [2:0] v_7332_0;
  reg [2:0] v_7333_0 = 3'h0;
  wire [0:0] v_7334_0;
  wire [0:0] v_7335_0;
  wire [0:0] v_7336_0;
  wire [2:0] v_7337_0;
  wire [2:0] v_7338_0;
  wire [2:0] v_7339_0;
  reg [2:0] v_7340_0 = 3'h0;
  wire [0:0] v_7341_0;
  wire [0:0] v_7342_0;
  wire [0:0] v_7343_0;
  wire [2:0] v_7344_0;
  wire [2:0] v_7345_0;
  wire [2:0] v_7346_0;
  reg [2:0] v_7347_0 = 3'h0;
  wire [0:0] v_7348_0;
  wire [0:0] v_7349_0;
  wire [0:0] v_7350_0;
  wire [2:0] v_7351_0;
  wire [2:0] v_7352_0;
  wire [2:0] v_7353_0;
  reg [2:0] v_7354_0 = 3'h0;
  wire [0:0] v_7355_0;
  wire [0:0] v_7356_0;
  wire [0:0] v_7357_0;
  wire [2:0] v_7358_0;
  wire [2:0] v_7359_0;
  wire [2:0] v_7360_0;
  reg [2:0] v_7361_0 = 3'h0;
  wire [0:0] v_7362_0;
  wire [0:0] v_7363_0;
  wire [0:0] v_7364_0;
  wire [2:0] v_7365_0;
  wire [2:0] v_7366_0;
  wire [2:0] v_7367_0;
  reg [2:0] v_7368_0 = 3'h0;
  wire [0:0] v_7369_0;
  wire [0:0] v_7370_0;
  wire [0:0] v_7371_0;
  wire [2:0] v_7372_0;
  wire [2:0] v_7373_0;
  wire [2:0] v_7374_0;
  reg [2:0] v_7375_0 = 3'h0;
  wire [0:0] v_7376_0;
  wire [0:0] v_7377_0;
  wire [0:0] v_7378_0;
  wire [2:0] v_7379_0;
  wire [2:0] v_7380_0;
  wire [2:0] v_7381_0;
  reg [2:0] v_7382_0 = 3'h0;
  wire [0:0] v_7383_0;
  wire [0:0] v_7384_0;
  wire [0:0] v_7385_0;
  wire [2:0] v_7386_0;
  wire [2:0] v_7387_0;
  wire [2:0] v_7388_0;
  reg [2:0] v_7389_0 = 3'h0;
  wire [0:0] v_7390_0;
  wire [0:0] v_7391_0;
  wire [0:0] v_7392_0;
  wire [2:0] v_7393_0;
  wire [2:0] v_7394_0;
  wire [2:0] v_7395_0;
  reg [2:0] v_7396_0 = 3'h0;
  wire [0:0] v_7397_0;
  wire [0:0] v_7398_0;
  wire [0:0] v_7399_0;
  wire [2:0] v_7400_0;
  wire [2:0] v_7401_0;
  wire [2:0] v_7402_0;
  reg [2:0] v_7403_0 = 3'h0;
  wire [0:0] v_7404_0;
  wire [0:0] v_7405_0;
  wire [0:0] v_7406_0;
  wire [2:0] v_7407_0;
  wire [2:0] v_7408_0;
  wire [2:0] v_7409_0;
  reg [2:0] v_7410_0 = 3'h0;
  wire [0:0] v_7411_0;
  wire [0:0] v_7412_0;
  wire [0:0] v_7413_0;
  wire [2:0] v_7414_0;
  wire [2:0] v_7415_0;
  wire [2:0] v_7416_0;
  reg [2:0] v_7417_0 = 3'h0;
  wire [0:0] v_7418_0;
  wire [0:0] v_7419_0;
  wire [0:0] v_7420_0;
  wire [2:0] v_7421_0;
  wire [2:0] v_7422_0;
  wire [2:0] v_7423_0;
  reg [2:0] v_7424_0 = 3'h0;
  wire [0:0] v_7425_0;
  wire [0:0] v_7426_0;
  wire [0:0] v_7427_0;
  wire [2:0] v_7428_0;
  wire [2:0] v_7429_0;
  wire [2:0] v_7430_0;
  reg [2:0] v_7431_0 = 3'h0;
  wire [0:0] v_7432_0;
  wire [0:0] v_7433_0;
  wire [0:0] v_7434_0;
  wire [2:0] v_7435_0;
  wire [2:0] v_7436_0;
  wire [2:0] v_7437_0;
  reg [2:0] v_7438_0 = 3'h0;
  wire [0:0] v_7439_0;
  wire [0:0] v_7440_0;
  wire [0:0] v_7441_0;
  wire [2:0] v_7442_0;
  wire [2:0] v_7443_0;
  wire [2:0] v_7444_0;
  reg [2:0] v_7445_0 = 3'h0;
  wire [0:0] v_7446_0;
  wire [0:0] v_7447_0;
  wire [0:0] v_7448_0;
  wire [2:0] v_7449_0;
  wire [2:0] v_7450_0;
  wire [2:0] v_7451_0;
  reg [2:0] v_7452_0 = 3'h0;
  wire [0:0] v_7453_0;
  wire [0:0] v_7454_0;
  wire [0:0] v_7455_0;
  wire [2:0] v_7456_0;
  wire [2:0] v_7457_0;
  wire [2:0] v_7458_0;
  reg [2:0] v_7459_0 = 3'h0;
  wire [0:0] v_7460_0;
  wire [0:0] v_7461_0;
  wire [0:0] v_7462_0;
  wire [2:0] v_7463_0;
  wire [2:0] v_7464_0;
  wire [2:0] v_7465_0;
  reg [2:0] v_7466_0 = 3'h0;
  wire [0:0] v_7467_0;
  wire [0:0] v_7468_0;
  wire [0:0] v_7469_0;
  wire [2:0] v_7470_0;
  wire [2:0] v_7471_0;
  wire [2:0] v_7472_0;
  reg [2:0] v_7473_0 = 3'h0;
  wire [0:0] v_7474_0;
  wire [0:0] v_7475_0;
  wire [0:0] v_7476_0;
  wire [2:0] v_7477_0;
  wire [2:0] v_7478_0;
  wire [2:0] v_7479_0;
  reg [2:0] v_7480_0 = 3'h0;
  wire [0:0] v_7481_0;
  wire [0:0] v_7482_0;
  wire [0:0] v_7483_0;
  wire [2:0] v_7484_0;
  wire [2:0] v_7485_0;
  wire [2:0] v_7486_0;
  reg [2:0] v_7487_0 = 3'h0;
  wire [0:0] v_7488_0;
  wire [0:0] v_7489_0;
  wire [0:0] v_7490_0;
  wire [2:0] v_7491_0;
  wire [2:0] v_7492_0;
  wire [2:0] v_7493_0;
  reg [2:0] v_7494_0 = 3'h0;
  wire [0:0] v_7495_0;
  wire [0:0] v_7496_0;
  wire [0:0] v_7497_0;
  wire [2:0] v_7498_0;
  wire [2:0] v_7499_0;
  wire [2:0] v_7500_0;
  reg [2:0] v_7501_0 = 3'h0;
  wire [0:0] v_7502_0;
  wire [0:0] v_7503_0;
  wire [0:0] v_7504_0;
  wire [2:0] v_7505_0;
  wire [2:0] v_7506_0;
  wire [2:0] v_7507_0;
  reg [2:0] v_7508_0 = 3'h0;
  wire [0:0] v_7509_0;
  wire [0:0] v_7510_0;
  wire [0:0] v_7511_0;
  wire [2:0] v_7512_0;
  wire [2:0] v_7513_0;
  wire [2:0] v_7514_0;
  reg [2:0] v_7515_0 = 3'h0;
  wire [0:0] v_7516_0;
  wire [0:0] v_7517_0;
  wire [0:0] v_7518_0;
  wire [2:0] v_7519_0;
  wire [2:0] v_7520_0;
  wire [2:0] v_7521_0;
  reg [2:0] v_7522_0 = 3'h0;
  wire [0:0] v_7523_0;
  wire [0:0] v_7524_0;
  wire [0:0] v_7525_0;
  wire [2:0] v_7526_0;
  wire [2:0] v_7527_0;
  wire [2:0] v_7528_0;
  reg [2:0] v_7529_0 = 3'h0;
  wire [0:0] v_7530_0;
  wire [0:0] v_7531_0;
  wire [0:0] v_7532_0;
  wire [2:0] v_7533_0;
  wire [2:0] v_7534_0;
  wire [2:0] v_7535_0;
  reg [2:0] v_7536_0 = 3'h0;
  wire [0:0] v_7537_0;
  wire [0:0] v_7538_0;
  wire [0:0] v_7539_0;
  wire [2:0] v_7540_0;
  wire [2:0] v_7541_0;
  wire [2:0] v_7542_0;
  reg [2:0] v_7543_0 = 3'h0;
  wire [0:0] v_7544_0;
  wire [0:0] v_7545_0;
  wire [0:0] v_7546_0;
  wire [2:0] v_7547_0;
  wire [2:0] v_7548_0;
  wire [2:0] v_7549_0;
  reg [2:0] v_7550_0 = 3'h0;
  wire [0:0] v_7551_0;
  wire [0:0] v_7552_0;
  wire [0:0] v_7553_0;
  wire [2:0] v_7554_0;
  wire [2:0] v_7555_0;
  wire [2:0] v_7556_0;
  reg [2:0] v_7557_0 = 3'h0;
  wire [0:0] v_7558_0;
  wire [0:0] v_7559_0;
  wire [0:0] v_7560_0;
  wire [2:0] v_7561_0;
  wire [2:0] v_7562_0;
  wire [2:0] v_7563_0;
  reg [2:0] v_7564_0 = 3'h0;
  wire [0:0] v_7565_0;
  wire [0:0] v_7566_0;
  wire [0:0] v_7567_0;
  wire [2:0] v_7568_0;
  wire [2:0] v_7569_0;
  wire [2:0] v_7570_0;
  reg [2:0] v_7571_0 = 3'h0;
  wire [0:0] v_7572_0;
  wire [0:0] v_7573_0;
  wire [0:0] v_7574_0;
  wire [2:0] v_7575_0;
  wire [2:0] v_7576_0;
  wire [2:0] v_7577_0;
  reg [2:0] v_7578_0 = 3'h0;
  wire [0:0] v_7579_0;
  wire [0:0] v_7580_0;
  wire [0:0] v_7581_0;
  wire [2:0] v_7582_0;
  wire [2:0] v_7583_0;
  wire [2:0] v_7584_0;
  reg [2:0] v_7585_0 = 3'h0;
  wire [0:0] v_7586_0;
  wire [0:0] v_7587_0;
  wire [0:0] v_7588_0;
  wire [2:0] v_7589_0;
  wire [2:0] v_7590_0;
  wire [2:0] v_7591_0;
  reg [2:0] v_7592_0 = 3'h0;
  wire [0:0] v_7593_0;
  wire [0:0] v_7594_0;
  wire [0:0] v_7595_0;
  wire [2:0] v_7596_0;
  wire [2:0] v_7597_0;
  wire [2:0] v_7598_0;
  reg [2:0] v_7599_0 = 3'h0;
  wire [0:0] v_7600_0;
  wire [0:0] v_7601_0;
  wire [0:0] v_7602_0;
  wire [2:0] v_7603_0;
  wire [2:0] v_7604_0;
  wire [2:0] v_7605_0;
  reg [2:0] v_7606_0 = 3'h0;
  wire [0:0] v_7607_0;
  wire [0:0] v_7608_0;
  wire [0:0] v_7609_0;
  wire [2:0] v_7610_0;
  wire [2:0] v_7611_0;
  wire [2:0] v_7612_0;
  reg [2:0] v_7613_0 = 3'h0;
  wire [0:0] v_7614_0;
  wire [0:0] v_7615_0;
  wire [0:0] v_7616_0;
  wire [2:0] v_7617_0;
  wire [2:0] v_7618_0;
  wire [2:0] v_7619_0;
  reg [2:0] v_7620_0 = 3'h0;
  wire [0:0] v_7621_0;
  wire [0:0] v_7622_0;
  wire [0:0] v_7623_0;
  wire [2:0] v_7624_0;
  wire [2:0] v_7625_0;
  wire [2:0] v_7626_0;
  reg [2:0] v_7627_0 = 3'h0;
  wire [0:0] v_7628_0;
  wire [0:0] v_7629_0;
  wire [0:0] v_7630_0;
  wire [2:0] v_7631_0;
  wire [2:0] v_7632_0;
  wire [2:0] v_7633_0;
  reg [2:0] v_7634_0 = 3'h0;
  wire [0:0] v_7635_0;
  wire [0:0] v_7636_0;
  wire [0:0] v_7637_0;
  wire [2:0] v_7638_0;
  wire [2:0] v_7639_0;
  wire [2:0] v_7640_0;
  reg [2:0] v_7641_0 = 3'h0;
  wire [0:0] v_7642_0;
  wire [0:0] v_7643_0;
  wire [0:0] v_7644_0;
  wire [2:0] v_7645_0;
  wire [2:0] v_7646_0;
  wire [2:0] v_7647_0;
  reg [2:0] v_7648_0 = 3'h0;
  wire [0:0] v_7649_0;
  wire [0:0] v_7650_0;
  wire [0:0] v_7651_0;
  wire [2:0] v_7652_0;
  wire [2:0] v_7653_0;
  wire [2:0] v_7654_0;
  reg [2:0] v_7655_0 = 3'h0;
  wire [0:0] v_7656_0;
  wire [0:0] v_7657_0;
  wire [0:0] v_7658_0;
  wire [2:0] v_7659_0;
  wire [2:0] v_7660_0;
  wire [2:0] v_7661_0;
  reg [2:0] v_7662_0 = 3'h0;
  wire [0:0] v_7663_0;
  wire [0:0] v_7664_0;
  wire [0:0] v_7665_0;
  wire [2:0] v_7666_0;
  wire [2:0] v_7667_0;
  wire [2:0] v_7668_0;
  reg [2:0] v_7669_0 = 3'h0;
  wire [0:0] v_7670_0;
  wire [0:0] v_7671_0;
  wire [0:0] v_7672_0;
  wire [2:0] v_7673_0;
  wire [2:0] v_7674_0;
  wire [2:0] v_7675_0;
  reg [2:0] v_7676_0 = 3'h0;
  wire [0:0] v_7677_0;
  wire [0:0] v_7678_0;
  wire [0:0] v_7679_0;
  wire [2:0] v_7680_0;
  wire [2:0] v_7681_0;
  wire [2:0] v_7682_0;
  reg [2:0] v_7683_0 = 3'h0;
  wire [0:0] v_7684_0;
  wire [0:0] v_7685_0;
  wire [0:0] v_7686_0;
  wire [2:0] v_7687_0;
  wire [2:0] v_7688_0;
  wire [2:0] v_7689_0;
  reg [2:0] v_7690_0 = 3'h0;
  wire [0:0] v_7691_0;
  wire [0:0] v_7692_0;
  wire [0:0] v_7693_0;
  wire [2:0] v_7694_0;
  wire [2:0] v_7695_0;
  wire [2:0] v_7696_0;
  reg [2:0] v_7697_0 = 3'h0;
  wire [0:0] v_7698_0;
  wire [0:0] v_7699_0;
  wire [0:0] v_7700_0;
  wire [2:0] v_7701_0;
  wire [2:0] v_7702_0;
  wire [2:0] v_7703_0;
  reg [2:0] v_7704_0 = 3'h0;
  wire [0:0] v_7705_0;
  wire [0:0] v_7706_0;
  wire [0:0] v_7707_0;
  wire [2:0] v_7708_0;
  wire [2:0] v_7709_0;
  wire [2:0] v_7710_0;
  reg [2:0] v_7711_0 = 3'h0;
  wire [0:0] v_7712_0;
  wire [0:0] v_7713_0;
  wire [0:0] v_7714_0;
  wire [2:0] v_7715_0;
  wire [2:0] v_7716_0;
  wire [2:0] v_7717_0;
  reg [2:0] v_7718_0 = 3'h0;
  wire [0:0] v_7719_0;
  wire [0:0] v_7720_0;
  wire [0:0] v_7721_0;
  wire [2:0] v_7722_0;
  wire [2:0] v_7723_0;
  wire [2:0] v_7724_0;
  reg [2:0] v_7725_0 = 3'h0;
  wire [0:0] v_7726_0;
  wire [0:0] v_7727_0;
  wire [0:0] v_7728_0;
  wire [2:0] v_7729_0;
  wire [2:0] v_7730_0;
  wire [2:0] v_7731_0;
  reg [2:0] v_7732_0 = 3'h0;
  wire [0:0] v_7733_0;
  wire [0:0] v_7734_0;
  wire [0:0] v_7735_0;
  wire [2:0] v_7736_0;
  wire [2:0] v_7737_0;
  wire [2:0] v_7738_0;
  reg [2:0] v_7739_0 = 3'h0;
  wire [0:0] v_7740_0;
  wire [0:0] v_7741_0;
  wire [0:0] v_7742_0;
  wire [2:0] v_7743_0;
  wire [2:0] v_7744_0;
  wire [2:0] v_7745_0;
  reg [2:0] v_7746_0 = 3'h0;
  wire [0:0] v_7747_0;
  wire [0:0] v_7748_0;
  wire [0:0] v_7749_0;
  wire [2:0] v_7750_0;
  wire [2:0] v_7751_0;
  wire [2:0] v_7752_0;
  reg [2:0] v_7753_0 = 3'h0;
  wire [0:0] v_7754_0;
  wire [0:0] v_7755_0;
  wire [0:0] v_7756_0;
  wire [2:0] v_7757_0;
  wire [2:0] v_7758_0;
  wire [2:0] v_7759_0;
  reg [2:0] v_7760_0 = 3'h0;
  wire [0:0] v_7761_0;
  wire [0:0] v_7762_0;
  wire [0:0] v_7763_0;
  wire [2:0] v_7764_0;
  wire [2:0] v_7765_0;
  wire [2:0] v_7766_0;
  reg [2:0] v_7767_0 = 3'h0;
  wire [0:0] v_7768_0;
  wire [0:0] v_7769_0;
  wire [0:0] v_7770_0;
  wire [2:0] v_7771_0;
  wire [2:0] v_7772_0;
  wire [2:0] v_7773_0;
  reg [2:0] v_7774_0 = 3'h0;
  wire [0:0] v_7775_0;
  wire [0:0] v_7776_0;
  wire [0:0] v_7777_0;
  wire [2:0] v_7778_0;
  wire [2:0] v_7779_0;
  wire [2:0] v_7780_0;
  reg [2:0] v_7781_0 = 3'h0;
  wire [0:0] v_7782_0;
  wire [0:0] v_7783_0;
  wire [0:0] v_7784_0;
  wire [2:0] v_7785_0;
  wire [2:0] v_7786_0;
  wire [2:0] v_7787_0;
  reg [2:0] v_7788_0 = 3'h0;
  wire [0:0] v_7789_0;
  wire [0:0] v_7790_0;
  wire [0:0] v_7791_0;
  wire [2:0] v_7792_0;
  wire [2:0] v_7793_0;
  wire [2:0] v_7794_0;
  reg [2:0] v_7795_0 = 3'h0;
  wire [0:0] v_7796_0;
  wire [0:0] v_7797_0;
  wire [0:0] v_7798_0;
  wire [2:0] v_7799_0;
  wire [2:0] v_7800_0;
  wire [2:0] v_7801_0;
  reg [2:0] v_7802_0 = 3'h0;
  wire [0:0] v_7803_0;
  wire [0:0] v_7804_0;
  wire [0:0] v_7805_0;
  wire [2:0] v_7806_0;
  wire [2:0] v_7807_0;
  wire [2:0] v_7808_0;
  reg [2:0] v_7809_0 = 3'h0;
  wire [0:0] v_7810_0;
  wire [0:0] v_7811_0;
  wire [0:0] v_7812_0;
  wire [2:0] v_7813_0;
  wire [2:0] v_7814_0;
  wire [2:0] v_7815_0;
  reg [2:0] v_7816_0 = 3'h0;
  wire [0:0] v_7817_0;
  wire [0:0] v_7818_0;
  wire [0:0] v_7819_0;
  wire [2:0] v_7820_0;
  wire [2:0] v_7821_0;
  wire [2:0] v_7822_0;
  reg [2:0] v_7823_0 = 3'h0;
  wire [0:0] v_7824_0;
  wire [0:0] v_7825_0;
  wire [0:0] v_7826_0;
  wire [2:0] v_7827_0;
  wire [2:0] v_7828_0;
  wire [2:0] v_7829_0;
  reg [2:0] v_7830_0 = 3'h0;
  wire [0:0] v_7831_0;
  wire [0:0] v_7832_0;
  wire [0:0] v_7833_0;
  wire [2:0] v_7834_0;
  wire [2:0] v_7835_0;
  wire [2:0] v_7836_0;
  reg [2:0] v_7837_0 = 3'h0;
  wire [0:0] v_7838_0;
  wire [0:0] v_7839_0;
  wire [0:0] v_7840_0;
  wire [2:0] v_7841_0;
  wire [2:0] v_7842_0;
  wire [2:0] v_7843_0;
  reg [2:0] v_7844_0 = 3'h0;
  wire [0:0] v_7845_0;
  wire [0:0] v_7846_0;
  wire [0:0] v_7847_0;
  wire [2:0] v_7848_0;
  wire [2:0] v_7849_0;
  wire [2:0] v_7850_0;
  reg [2:0] v_7851_0 = 3'h0;
  wire [0:0] v_7852_0;
  wire [2:0] v_7853_0;
  wire [2:0] v_7854_0;
  wire [2:0] v_7855_0;
  wire [2:0] v_7856_0;
  wire [2:0] v_7857_0;
  wire [2:0] v_7858_0;
  wire [2:0] v_7859_0;
  wire [2:0] v_7860_0;
  wire [2:0] v_7861_0;
  wire [2:0] v_7862_0;
  wire [2:0] v_7863_0;
  wire [2:0] v_7864_0;
  wire [2:0] v_7865_0;
  wire [2:0] v_7866_0;
  wire [2:0] v_7867_0;
  wire [2:0] v_7868_0;
  wire [2:0] v_7869_0;
  wire [2:0] v_7870_0;
  wire [2:0] v_7871_0;
  wire [2:0] v_7872_0;
  wire [2:0] v_7873_0;
  wire [2:0] v_7874_0;
  wire [2:0] v_7875_0;
  wire [2:0] v_7876_0;
  wire [2:0] v_7877_0;
  wire [2:0] v_7878_0;
  wire [2:0] v_7879_0;
  wire [2:0] v_7880_0;
  wire [2:0] v_7881_0;
  wire [2:0] v_7882_0;
  wire [2:0] v_7883_0;
  wire [2:0] v_7884_0;
  wire [2:0] v_7885_0;
  wire [2:0] v_7886_0;
  wire [2:0] v_7887_0;
  wire [2:0] v_7888_0;
  wire [2:0] v_7889_0;
  wire [2:0] v_7890_0;
  wire [2:0] v_7891_0;
  wire [2:0] v_7892_0;
  wire [2:0] v_7893_0;
  wire [2:0] v_7894_0;
  wire [2:0] v_7895_0;
  wire [2:0] v_7896_0;
  wire [2:0] v_7897_0;
  wire [2:0] v_7898_0;
  wire [2:0] v_7899_0;
  wire [2:0] v_7900_0;
  wire [2:0] v_7901_0;
  wire [2:0] v_7902_0;
  wire [2:0] v_7903_0;
  wire [2:0] v_7904_0;
  wire [2:0] v_7905_0;
  wire [2:0] v_7906_0;
  wire [2:0] v_7907_0;
  wire [2:0] v_7908_0;
  wire [2:0] v_7909_0;
  wire [2:0] v_7910_0;
  wire [2:0] v_7911_0;
  wire [2:0] v_7912_0;
  wire [2:0] v_7913_0;
  wire [2:0] v_7914_0;
  wire [2:0] v_7915_0;
  wire [2:0] v_7916_0;
  wire [2:0] v_7917_0;
  wire [2:0] v_7918_0;
  wire [2:0] v_7919_0;
  wire [2:0] v_7920_0;
  wire [2:0] v_7921_0;
  wire [2:0] v_7922_0;
  wire [2:0] v_7923_0;
  wire [2:0] v_7924_0;
  wire [2:0] v_7925_0;
  wire [2:0] v_7926_0;
  wire [2:0] v_7927_0;
  wire [2:0] v_7928_0;
  wire [2:0] v_7929_0;
  wire [2:0] v_7930_0;
  wire [2:0] v_7931_0;
  wire [2:0] v_7932_0;
  wire [2:0] v_7933_0;
  wire [2:0] v_7934_0;
  wire [2:0] v_7935_0;
  wire [2:0] v_7936_0;
  wire [2:0] v_7937_0;
  wire [2:0] v_7938_0;
  wire [2:0] v_7939_0;
  wire [2:0] v_7940_0;
  wire [2:0] v_7941_0;
  wire [2:0] v_7942_0;
  wire [2:0] v_7943_0;
  wire [2:0] v_7944_0;
  wire [2:0] v_7945_0;
  wire [2:0] v_7946_0;
  wire [2:0] v_7947_0;
  wire [2:0] v_7948_0;
  wire [2:0] v_7949_0;
  wire [2:0] v_7950_0;
  wire [2:0] v_7951_0;
  wire [2:0] v_7952_0;
  wire [2:0] v_7953_0;
  wire [2:0] v_7954_0;
  wire [2:0] v_7955_0;
  wire [2:0] v_7956_0;
  wire [2:0] v_7957_0;
  wire [2:0] v_7958_0;
  wire [2:0] v_7959_0;
  wire [2:0] v_7960_0;
  wire [2:0] v_7961_0;
  wire [2:0] v_7962_0;
  wire [2:0] v_7963_0;
  wire [2:0] v_7964_0;
  wire [2:0] v_7965_0;
  wire [2:0] v_7966_0;
  wire [2:0] v_7967_0;
  wire [2:0] v_7968_0;
  wire [2:0] v_7969_0;
  wire [2:0] v_7970_0;
  wire [2:0] v_7971_0;
  wire [2:0] v_7972_0;
  wire [2:0] v_7973_0;
  wire [2:0] v_7974_0;
  wire [2:0] v_7975_0;
  wire [2:0] v_7976_0;
  wire [2:0] v_7977_0;
  wire [2:0] v_7978_0;
  wire [2:0] v_7979_0;
  wire [2:0] v_7980_0;
  wire [2:0] v_7981_0;
  wire [2:0] v_7982_0;
  wire [2:0] v_7983_0;
  wire [2:0] v_7984_0;
  wire [2:0] v_7985_0;
  wire [2:0] v_7986_0;
  wire [2:0] v_7987_0;
  wire [2:0] v_7988_0;
  wire [2:0] v_7989_0;
  wire [2:0] v_7990_0;
  wire [2:0] v_7991_0;
  wire [2:0] v_7992_0;
  wire [2:0] v_7993_0;
  wire [2:0] v_7994_0;
  wire [2:0] v_7995_0;
  wire [2:0] v_7996_0;
  wire [2:0] v_7997_0;
  wire [2:0] v_7998_0;
  wire [2:0] v_7999_0;
  wire [2:0] v_8000_0;
  wire [2:0] v_8001_0;
  wire [2:0] v_8002_0;
  wire [2:0] v_8003_0;
  wire [2:0] v_8004_0;
  wire [2:0] v_8005_0;
  wire [2:0] v_8006_0;
  wire [2:0] v_8007_0;
  wire [2:0] v_8008_0;
  wire [2:0] v_8009_0;
  wire [2:0] v_8010_0;
  wire [2:0] v_8011_0;
  wire [2:0] v_8012_0;
  wire [2:0] v_8013_0;
  wire [2:0] v_8014_0;
  wire [2:0] v_8015_0;
  wire [2:0] v_8016_0;
  wire [2:0] v_8017_0;
  wire [2:0] v_8018_0;
  wire [2:0] v_8019_0;
  wire [2:0] v_8020_0;
  wire [2:0] v_8021_0;
  wire [2:0] v_8022_0;
  wire [2:0] v_8023_0;
  wire [2:0] v_8024_0;
  wire [2:0] v_8025_0;
  wire [2:0] v_8026_0;
  wire [2:0] v_8027_0;
  wire [2:0] v_8028_0;
  wire [2:0] v_8029_0;
  wire [2:0] v_8030_0;
  wire [2:0] v_8031_0;
  wire [2:0] v_8032_0;
  wire [2:0] v_8033_0;
  wire [2:0] v_8034_0;
  wire [2:0] v_8035_0;
  wire [2:0] v_8036_0;
  wire [2:0] v_8037_0;
  wire [2:0] v_8038_0;
  wire [2:0] v_8039_0;
  wire [2:0] v_8040_0;
  wire [2:0] v_8041_0;
  wire [2:0] v_8042_0;
  wire [2:0] v_8043_0;
  wire [2:0] v_8044_0;
  wire [2:0] v_8045_0;
  wire [2:0] v_8046_0;
  wire [2:0] v_8047_0;
  wire [2:0] v_8048_0;
  wire [2:0] v_8049_0;
  wire [2:0] v_8050_0;
  wire [2:0] v_8051_0;
  wire [2:0] v_8052_0;
  wire [2:0] v_8053_0;
  wire [2:0] v_8054_0;
  wire [2:0] v_8055_0;
  wire [2:0] v_8056_0;
  wire [2:0] v_8057_0;
  wire [2:0] v_8058_0;
  wire [2:0] v_8059_0;
  wire [2:0] v_8060_0;
  wire [2:0] v_8061_0;
  wire [2:0] v_8062_0;
  wire [2:0] v_8063_0;
  wire [2:0] v_8064_0;
  wire [2:0] v_8065_0;
  wire [2:0] v_8066_0;
  wire [2:0] v_8067_0;
  wire [2:0] v_8068_0;
  wire [2:0] v_8069_0;
  wire [2:0] v_8070_0;
  wire [2:0] v_8071_0;
  wire [2:0] v_8072_0;
  wire [2:0] v_8073_0;
  wire [2:0] v_8074_0;
  wire [2:0] v_8075_0;
  wire [2:0] v_8076_0;
  wire [2:0] v_8077_0;
  wire [2:0] v_8078_0;
  wire [2:0] v_8079_0;
  wire [2:0] v_8080_0;
  wire [2:0] v_8081_0;
  wire [2:0] v_8082_0;
  wire [2:0] v_8083_0;
  wire [2:0] v_8084_0;
  wire [2:0] v_8085_0;
  wire [2:0] v_8086_0;
  wire [2:0] v_8087_0;
  wire [2:0] v_8088_0;
  wire [2:0] v_8089_0;
  wire [2:0] v_8090_0;
  wire [2:0] v_8091_0;
  wire [2:0] v_8092_0;
  wire [2:0] v_8093_0;
  wire [2:0] v_8094_0;
  wire [2:0] v_8095_0;
  wire [2:0] v_8096_0;
  wire [2:0] v_8097_0;
  wire [2:0] v_8098_0;
  wire [2:0] v_8099_0;
  wire [2:0] v_8100_0;
  wire [2:0] v_8101_0;
  wire [2:0] v_8102_0;
  wire [2:0] v_8103_0;
  wire [2:0] v_8104_0;
  wire [2:0] v_8105_0;
  wire [2:0] v_8106_0;
  wire [2:0] v_8107_0;
  wire [2:0] v_8108_0;
  wire [2:0] v_8109_0;
  wire [2:0] v_8110_0;
  wire [2:0] v_8111_0;
  wire [2:0] v_8112_0;
  wire [2:0] v_8113_0;
  wire [2:0] v_8114_0;
  wire [2:0] v_8115_0;
  wire [2:0] v_8116_0;
  wire [2:0] v_8117_0;
  wire [2:0] v_8118_0;
  wire [2:0] v_8119_0;
  wire [2:0] v_8120_0;
  wire [2:0] v_8121_0;
  wire [2:0] v_8122_0;
  wire [2:0] v_8123_0;
  wire [2:0] v_8124_0;
  wire [2:0] v_8125_0;
  wire [2:0] v_8126_0;
  wire [2:0] v_8127_0;
  wire [2:0] v_8128_0;
  wire [2:0] v_8129_0;
  wire [2:0] v_8130_0;
  wire [2:0] v_8131_0;
  wire [2:0] v_8132_0;
  wire [2:0] v_8133_0;
  wire [2:0] v_8134_0;
  wire [2:0] v_8135_0;
  wire [2:0] v_8136_0;
  wire [2:0] v_8137_0;
  wire [2:0] v_8138_0;
  wire [2:0] v_8139_0;
  wire [2:0] v_8140_0;
  wire [2:0] v_8141_0;
  wire [2:0] v_8142_0;
  wire [2:0] v_8143_0;
  wire [2:0] v_8144_0;
  wire [2:0] v_8145_0;
  wire [2:0] v_8146_0;
  wire [2:0] v_8147_0;
  wire [2:0] v_8148_0;
  wire [2:0] v_8149_0;
  wire [2:0] v_8150_0;
  wire [2:0] v_8151_0;
  wire [2:0] v_8152_0;
  wire [2:0] v_8153_0;
  wire [2:0] v_8154_0;
  wire [2:0] v_8155_0;
  wire [2:0] v_8156_0;
  wire [2:0] v_8157_0;
  wire [2:0] v_8158_0;
  wire [2:0] v_8159_0;
  wire [2:0] v_8160_0;
  wire [2:0] v_8161_0;
  wire [2:0] v_8162_0;
  wire [2:0] v_8163_0;
  wire [2:0] v_8164_0;
  wire [2:0] v_8165_0;
  wire [2:0] v_8166_0;
  wire [2:0] v_8167_0;
  wire [2:0] v_8168_0;
  wire [2:0] v_8169_0;
  wire [2:0] v_8170_0;
  wire [2:0] v_8171_0;
  wire [2:0] v_8172_0;
  wire [2:0] v_8173_0;
  wire [2:0] v_8174_0;
  wire [2:0] v_8175_0;
  wire [2:0] v_8176_0;
  wire [2:0] v_8177_0;
  wire [2:0] v_8178_0;
  wire [2:0] v_8179_0;
  wire [2:0] v_8180_0;
  wire [2:0] v_8181_0;
  wire [2:0] v_8182_0;
  wire [2:0] v_8183_0;
  wire [2:0] v_8184_0;
  wire [2:0] v_8185_0;
  wire [2:0] v_8186_0;
  wire [2:0] v_8187_0;
  wire [2:0] v_8188_0;
  wire [2:0] v_8189_0;
  wire [2:0] v_8190_0;
  wire [2:0] v_8191_0;
  wire [2:0] v_8192_0;
  wire [2:0] v_8193_0;
  wire [2:0] v_8194_0;
  wire [2:0] v_8195_0;
  wire [2:0] v_8196_0;
  wire [2:0] v_8197_0;
  wire [2:0] v_8198_0;
  wire [2:0] v_8199_0;
  wire [2:0] v_8200_0;
  wire [2:0] v_8201_0;
  wire [2:0] v_8202_0;
  wire [2:0] v_8203_0;
  wire [2:0] v_8204_0;
  wire [2:0] v_8205_0;
  wire [2:0] v_8206_0;
  wire [2:0] v_8207_0;
  wire [2:0] v_8208_0;
  wire [2:0] v_8209_0;
  wire [2:0] v_8210_0;
  wire [2:0] v_8211_0;
  wire [2:0] v_8212_0;
  wire [2:0] v_8213_0;
  wire [2:0] v_8214_0;
  wire [2:0] v_8215_0;
  wire [2:0] v_8216_0;
  wire [2:0] v_8217_0;
  wire [2:0] v_8218_0;
  wire [2:0] v_8219_0;
  wire [2:0] v_8220_0;
  wire [2:0] v_8221_0;
  wire [2:0] v_8222_0;
  wire [2:0] v_8223_0;
  wire [2:0] v_8224_0;
  wire [2:0] v_8225_0;
  wire [2:0] v_8226_0;
  wire [2:0] v_8227_0;
  wire [2:0] v_8228_0;
  wire [2:0] v_8229_0;
  wire [2:0] v_8230_0;
  wire [2:0] v_8231_0;
  wire [2:0] v_8232_0;
  wire [2:0] v_8233_0;
  wire [2:0] v_8234_0;
  wire [2:0] v_8235_0;
  wire [2:0] v_8236_0;
  wire [2:0] v_8237_0;
  wire [2:0] v_8238_0;
  wire [2:0] v_8239_0;
  wire [2:0] v_8240_0;
  wire [2:0] v_8241_0;
  wire [2:0] v_8242_0;
  wire [2:0] v_8243_0;
  wire [2:0] v_8244_0;
  wire [2:0] v_8245_0;
  wire [2:0] v_8246_0;
  wire [2:0] v_8247_0;
  wire [2:0] v_8248_0;
  wire [2:0] v_8249_0;
  wire [2:0] v_8250_0;
  wire [2:0] v_8251_0;
  wire [2:0] v_8252_0;
  wire [2:0] v_8253_0;
  wire [2:0] v_8254_0;
  wire [2:0] v_8255_0;
  wire [2:0] v_8256_0;
  wire [2:0] v_8257_0;
  wire [2:0] v_8258_0;
  wire [2:0] v_8259_0;
  wire [2:0] v_8260_0;
  wire [2:0] v_8261_0;
  wire [2:0] v_8262_0;
  wire [2:0] v_8263_0;
  wire [2:0] v_8264_0;
  wire [2:0] v_8265_0;
  wire [2:0] v_8266_0;
  wire [2:0] v_8267_0;
  wire [2:0] v_8268_0;
  wire [2:0] v_8269_0;
  wire [2:0] v_8270_0;
  wire [2:0] v_8271_0;
  wire [2:0] v_8272_0;
  wire [2:0] v_8273_0;
  wire [2:0] v_8274_0;
  wire [2:0] v_8275_0;
  wire [2:0] v_8276_0;
  wire [2:0] v_8277_0;
  wire [2:0] v_8278_0;
  wire [2:0] v_8279_0;
  wire [2:0] v_8280_0;
  wire [2:0] v_8281_0;
  wire [2:0] v_8282_0;
  wire [2:0] v_8283_0;
  wire [2:0] v_8284_0;
  wire [2:0] v_8285_0;
  wire [2:0] v_8286_0;
  wire [2:0] v_8287_0;
  wire [2:0] v_8288_0;
  wire [2:0] v_8289_0;
  wire [2:0] v_8290_0;
  wire [2:0] v_8291_0;
  wire [2:0] v_8292_0;
  wire [2:0] v_8293_0;
  wire [2:0] v_8294_0;
  wire [2:0] v_8295_0;
  wire [2:0] v_8296_0;
  wire [2:0] v_8297_0;
  wire [2:0] v_8298_0;
  wire [2:0] v_8299_0;
  wire [2:0] v_8300_0;
  wire [2:0] v_8301_0;
  wire [2:0] v_8302_0;
  wire [2:0] v_8303_0;
  wire [2:0] v_8304_0;
  wire [2:0] v_8305_0;
  wire [2:0] v_8306_0;
  wire [2:0] v_8307_0;
  wire [2:0] v_8308_0;
  wire [2:0] v_8309_0;
  wire [2:0] v_8310_0;
  wire [2:0] v_8311_0;
  wire [2:0] v_8312_0;
  wire [2:0] v_8313_0;
  wire [2:0] v_8314_0;
  wire [2:0] v_8315_0;
  wire [2:0] v_8316_0;
  wire [2:0] v_8317_0;
  wire [2:0] v_8318_0;
  wire [2:0] v_8319_0;
  wire [2:0] v_8320_0;
  wire [2:0] v_8321_0;
  wire [2:0] v_8322_0;
  wire [2:0] v_8323_0;
  wire [2:0] v_8324_0;
  wire [2:0] v_8325_0;
  wire [2:0] v_8326_0;
  wire [2:0] v_8327_0;
  wire [2:0] v_8328_0;
  wire [2:0] v_8329_0;
  wire [2:0] v_8330_0;
  wire [2:0] v_8331_0;
  wire [2:0] v_8332_0;
  wire [2:0] v_8333_0;
  wire [2:0] v_8334_0;
  wire [2:0] v_8335_0;
  wire [2:0] v_8336_0;
  wire [2:0] v_8337_0;
  wire [2:0] v_8338_0;
  wire [2:0] v_8339_0;
  wire [2:0] v_8340_0;
  wire [2:0] v_8341_0;
  wire [2:0] v_8342_0;
  wire [2:0] v_8343_0;
  wire [2:0] v_8344_0;
  wire [2:0] v_8345_0;
  wire [2:0] v_8346_0;
  wire [2:0] v_8347_0;
  wire [2:0] v_8348_0;
  wire [2:0] v_8349_0;
  wire [2:0] v_8350_0;
  wire [2:0] v_8351_0;
  wire [2:0] v_8352_0;
  wire [2:0] v_8353_0;
  wire [2:0] v_8354_0;
  wire [2:0] v_8355_0;
  wire [2:0] v_8356_0;
  wire [2:0] v_8357_0;
  wire [2:0] v_8358_0;
  wire [2:0] v_8359_0;
  wire [2:0] v_8360_0;
  wire [2:0] v_8361_0;
  wire [2:0] v_8362_0;
  wire [2:0] v_8363_0;
  wire [2:0] v_8364_0;
  wire [2:0] v_8365_0;
  wire [2:0] v_8366_0;
  wire [2:0] v_8367_0;
  wire [2:0] v_8368_0;
  wire [2:0] v_8369_0;
  wire [2:0] v_8370_0;
  wire [2:0] v_8371_0;
  wire [2:0] v_8372_0;
  wire [2:0] v_8373_0;
  wire [2:0] v_8374_0;
  wire [2:0] v_8375_0;
  wire [2:0] v_8376_0;
  wire [2:0] v_8377_0;
  wire [2:0] v_8378_0;
  wire [2:0] v_8379_0;
  wire [2:0] v_8380_0;
  wire [2:0] v_8381_0;
  wire [2:0] v_8382_0;
  wire [2:0] v_8383_0;
  wire [2:0] v_8384_0;
  wire [2:0] v_8385_0;
  wire [2:0] v_8386_0;
  wire [2:0] v_8387_0;
  wire [2:0] v_8388_0;
  wire [2:0] v_8389_0;
  wire [2:0] v_8390_0;
  wire [2:0] v_8391_0;
  wire [2:0] v_8392_0;
  wire [2:0] v_8393_0;
  wire [2:0] v_8394_0;
  wire [2:0] v_8395_0;
  wire [2:0] v_8396_0;
  wire [2:0] v_8397_0;
  wire [2:0] v_8398_0;
  wire [2:0] v_8399_0;
  wire [2:0] v_8400_0;
  wire [2:0] v_8401_0;
  wire [2:0] v_8402_0;
  wire [2:0] v_8403_0;
  wire [2:0] v_8404_0;
  wire [2:0] v_8405_0;
  wire [2:0] v_8406_0;
  wire [2:0] v_8407_0;
  wire [2:0] v_8408_0;
  wire [2:0] v_8409_0;
  wire [2:0] v_8410_0;
  wire [2:0] v_8411_0;
  wire [2:0] v_8412_0;
  wire [2:0] v_8413_0;
  wire [2:0] v_8414_0;
  wire [2:0] v_8415_0;
  wire [2:0] v_8416_0;
  wire [2:0] v_8417_0;
  wire [2:0] v_8418_0;
  wire [2:0] v_8419_0;
  wire [2:0] v_8420_0;
  wire [2:0] v_8421_0;
  wire [2:0] v_8422_0;
  wire [2:0] v_8423_0;
  wire [2:0] v_8424_0;
  wire [2:0] v_8425_0;
  wire [2:0] v_8426_0;
  wire [2:0] v_8427_0;
  wire [2:0] v_8428_0;
  wire [2:0] v_8429_0;
  wire [2:0] v_8430_0;
  wire [2:0] v_8431_0;
  wire [2:0] v_8432_0;
  wire [2:0] v_8433_0;
  wire [2:0] v_8434_0;
  wire [2:0] v_8435_0;
  wire [2:0] v_8436_0;
  wire [2:0] v_8437_0;
  wire [2:0] v_8438_0;
  wire [2:0] v_8439_0;
  wire [2:0] v_8440_0;
  wire [2:0] v_8441_0;
  wire [2:0] v_8442_0;
  wire [2:0] v_8443_0;
  wire [2:0] v_8444_0;
  wire [2:0] v_8445_0;
  wire [2:0] v_8446_0;
  wire [2:0] v_8447_0;
  wire [2:0] v_8448_0;
  wire [2:0] v_8449_0;
  wire [2:0] v_8450_0;
  wire [2:0] v_8451_0;
  wire [2:0] v_8452_0;
  wire [2:0] v_8453_0;
  wire [2:0] v_8454_0;
  wire [2:0] v_8455_0;
  wire [2:0] v_8456_0;
  wire [2:0] v_8457_0;
  wire [2:0] v_8458_0;
  wire [2:0] v_8459_0;
  wire [2:0] v_8460_0;
  wire [2:0] v_8461_0;
  wire [2:0] v_8462_0;
  wire [2:0] v_8463_0;
  wire [2:0] v_8464_0;
  wire [2:0] v_8465_0;
  wire [2:0] v_8466_0;
  wire [2:0] v_8467_0;
  wire [2:0] v_8468_0;
  wire [2:0] v_8469_0;
  wire [2:0] v_8470_0;
  wire [2:0] v_8471_0;
  wire [2:0] v_8472_0;
  wire [2:0] v_8473_0;
  wire [2:0] v_8474_0;
  wire [2:0] v_8475_0;
  wire [2:0] v_8476_0;
  wire [2:0] v_8477_0;
  wire [2:0] v_8478_0;
  wire [2:0] v_8479_0;
  wire [2:0] v_8480_0;
  wire [2:0] v_8481_0;
  wire [2:0] v_8482_0;
  wire [2:0] v_8483_0;
  wire [2:0] v_8484_0;
  wire [2:0] v_8485_0;
  wire [2:0] v_8486_0;
  wire [2:0] v_8487_0;
  wire [2:0] v_8488_0;
  wire [2:0] v_8489_0;
  wire [2:0] v_8490_0;
  wire [2:0] v_8491_0;
  wire [2:0] v_8492_0;
  wire [2:0] v_8493_0;
  wire [2:0] v_8494_0;
  wire [2:0] v_8495_0;
  wire [2:0] v_8496_0;
  wire [2:0] v_8497_0;
  wire [2:0] v_8498_0;
  wire [2:0] v_8499_0;
  wire [2:0] v_8500_0;
  wire [2:0] v_8501_0;
  wire [2:0] v_8502_0;
  wire [2:0] v_8503_0;
  wire [2:0] v_8504_0;
  wire [2:0] v_8505_0;
  wire [2:0] v_8506_0;
  wire [2:0] v_8507_0;
  wire [2:0] v_8508_0;
  wire [2:0] v_8509_0;
  wire [2:0] v_8510_0;
  wire [2:0] v_8511_0;
  wire [2:0] v_8512_0;
  wire [2:0] v_8513_0;
  wire [2:0] v_8514_0;
  wire [2:0] v_8515_0;
  wire [2:0] v_8516_0;
  wire [2:0] v_8517_0;
  wire [2:0] v_8518_0;
  wire [2:0] v_8519_0;
  wire [2:0] v_8520_0;
  wire [2:0] v_8521_0;
  wire [2:0] v_8522_0;
  wire [2:0] v_8523_0;
  wire [2:0] v_8524_0;
  wire [2:0] v_8525_0;
  wire [2:0] v_8526_0;
  wire [2:0] v_8527_0;
  wire [2:0] v_8528_0;
  wire [2:0] v_8529_0;
  wire [2:0] v_8530_0;
  wire [2:0] v_8531_0;
  wire [2:0] v_8532_0;
  wire [2:0] v_8533_0;
  wire [2:0] v_8534_0;
  wire [2:0] v_8535_0;
  wire [2:0] v_8536_0;
  wire [2:0] v_8537_0;
  wire [2:0] v_8538_0;
  wire [2:0] v_8539_0;
  wire [2:0] v_8540_0;
  wire [2:0] v_8541_0;
  wire [2:0] v_8542_0;
  wire [2:0] v_8543_0;
  wire [2:0] v_8544_0;
  wire [2:0] v_8545_0;
  wire [2:0] v_8546_0;
  wire [2:0] v_8547_0;
  wire [2:0] v_8548_0;
  wire [2:0] v_8549_0;
  wire [2:0] v_8550_0;
  wire [2:0] v_8551_0;
  wire [2:0] v_8552_0;
  wire [2:0] v_8553_0;
  wire [2:0] v_8554_0;
  wire [2:0] v_8555_0;
  wire [2:0] v_8556_0;
  wire [2:0] v_8557_0;
  wire [2:0] v_8558_0;
  wire [2:0] v_8559_0;
  wire [2:0] v_8560_0;
  wire [2:0] v_8561_0;
  wire [2:0] v_8562_0;
  wire [2:0] v_8563_0;
  wire [2:0] v_8564_0;
  wire [2:0] v_8565_0;
  wire [2:0] v_8566_0;
  wire [2:0] v_8567_0;
  wire [2:0] v_8568_0;
  wire [2:0] v_8569_0;
  wire [2:0] v_8570_0;
  wire [2:0] v_8571_0;
  wire [2:0] v_8572_0;
  wire [2:0] v_8573_0;
  wire [2:0] v_8574_0;
  wire [2:0] v_8575_0;
  wire [2:0] v_8576_0;
  wire [2:0] v_8577_0;
  wire [2:0] v_8578_0;
  wire [2:0] v_8579_0;
  wire [2:0] v_8580_0;
  wire [2:0] v_8581_0;
  wire [2:0] v_8582_0;
  wire [2:0] v_8583_0;
  wire [2:0] v_8584_0;
  wire [2:0] v_8585_0;
  wire [2:0] v_8586_0;
  wire [2:0] v_8587_0;
  wire [2:0] v_8588_0;
  wire [2:0] v_8589_0;
  wire [2:0] v_8590_0;
  wire [2:0] v_8591_0;
  wire [2:0] v_8592_0;
  wire [2:0] v_8593_0;
  wire [2:0] v_8594_0;
  wire [2:0] v_8595_0;
  wire [2:0] v_8596_0;
  wire [2:0] v_8597_0;
  wire [2:0] v_8598_0;
  wire [2:0] v_8599_0;
  wire [2:0] v_8600_0;
  wire [2:0] v_8601_0;
  wire [2:0] v_8602_0;
  wire [2:0] v_8603_0;
  wire [2:0] v_8604_0;
  wire [2:0] v_8605_0;
  wire [2:0] v_8606_0;
  wire [2:0] v_8607_0;
  wire [2:0] v_8608_0;
  wire [2:0] v_8609_0;
  wire [2:0] v_8610_0;
  wire [2:0] v_8611_0;
  wire [2:0] v_8612_0;
  wire [2:0] v_8613_0;
  wire [2:0] v_8614_0;
  wire [2:0] v_8615_0;
  wire [2:0] v_8616_0;
  wire [2:0] v_8617_0;
  wire [2:0] v_8618_0;
  wire [2:0] v_8619_0;
  wire [2:0] v_8620_0;
  wire [2:0] v_8621_0;
  wire [2:0] v_8622_0;
  wire [2:0] v_8623_0;
  wire [2:0] v_8624_0;
  wire [2:0] v_8625_0;
  wire [2:0] v_8626_0;
  wire [2:0] v_8627_0;
  wire [2:0] v_8628_0;
  wire [2:0] v_8629_0;
  wire [2:0] v_8630_0;
  wire [2:0] v_8631_0;
  wire [2:0] v_8632_0;
  wire [2:0] v_8633_0;
  wire [2:0] v_8634_0;
  wire [2:0] v_8635_0;
  wire [2:0] v_8636_0;
  wire [2:0] v_8637_0;
  wire [2:0] v_8638_0;
  wire [2:0] v_8639_0;
  wire [2:0] v_8640_0;
  wire [2:0] v_8641_0;
  wire [2:0] v_8642_0;
  wire [2:0] v_8643_0;
  wire [2:0] v_8644_0;
  wire [2:0] v_8645_0;
  wire [2:0] v_8646_0;
  wire [2:0] v_8647_0;
  wire [2:0] v_8648_0;
  wire [2:0] v_8649_0;
  wire [2:0] v_8650_0;
  wire [2:0] v_8651_0;
  wire [2:0] v_8652_0;
  wire [2:0] v_8653_0;
  wire [2:0] v_8654_0;
  wire [2:0] v_8655_0;
  wire [2:0] v_8656_0;
  wire [2:0] v_8657_0;
  wire [2:0] v_8658_0;
  wire [2:0] v_8659_0;
  wire [2:0] v_8660_0;
  wire [2:0] v_8661_0;
  wire [2:0] v_8662_0;
  wire [2:0] v_8663_0;
  wire [2:0] v_8664_0;
  wire [2:0] v_8665_0;
  wire [2:0] v_8666_0;
  wire [2:0] v_8667_0;
  wire [2:0] v_8668_0;
  wire [2:0] v_8669_0;
  wire [2:0] v_8670_0;
  wire [2:0] v_8671_0;
  wire [2:0] v_8672_0;
  wire [2:0] v_8673_0;
  wire [2:0] v_8674_0;
  wire [2:0] v_8675_0;
  wire [2:0] v_8676_0;
  wire [2:0] v_8677_0;
  wire [2:0] v_8678_0;
  wire [2:0] v_8679_0;
  wire [2:0] v_8680_0;
  wire [2:0] v_8681_0;
  wire [2:0] v_8682_0;
  wire [2:0] v_8683_0;
  wire [2:0] v_8684_0;
  wire [2:0] v_8685_0;
  wire [2:0] v_8686_0;
  wire [2:0] v_8687_0;
  wire [2:0] v_8688_0;
  wire [2:0] v_8689_0;
  wire [2:0] v_8690_0;
  wire [2:0] v_8691_0;
  wire [2:0] v_8692_0;
  wire [2:0] v_8693_0;
  wire [2:0] v_8694_0;
  wire [2:0] v_8695_0;
  wire [2:0] v_8696_0;
  wire [2:0] v_8697_0;
  wire [2:0] v_8698_0;
  wire [2:0] v_8699_0;
  wire [2:0] v_8700_0;
  wire [2:0] v_8701_0;
  wire [2:0] v_8702_0;
  wire [2:0] v_8703_0;
  wire [2:0] v_8704_0;
  wire [2:0] v_8705_0;
  wire [2:0] v_8706_0;
  wire [2:0] v_8707_0;
  wire [2:0] v_8708_0;
  wire [2:0] v_8709_0;
  wire [2:0] v_8710_0;
  wire [2:0] v_8711_0;
  wire [2:0] v_8712_0;
  wire [2:0] v_8713_0;
  wire [2:0] v_8714_0;
  wire [2:0] v_8715_0;
  wire [2:0] v_8716_0;
  wire [2:0] v_8717_0;
  wire [2:0] v_8718_0;
  wire [2:0] v_8719_0;
  wire [2:0] v_8720_0;
  wire [2:0] v_8721_0;
  wire [2:0] v_8722_0;
  wire [2:0] v_8723_0;
  wire [2:0] v_8724_0;
  wire [2:0] v_8725_0;
  wire [2:0] v_8726_0;
  wire [2:0] v_8727_0;
  wire [2:0] v_8728_0;
  wire [2:0] v_8729_0;
  wire [2:0] v_8730_0;
  wire [2:0] v_8731_0;
  wire [2:0] v_8732_0;
  wire [2:0] v_8733_0;
  wire [2:0] v_8734_0;
  wire [2:0] v_8735_0;
  wire [2:0] v_8736_0;
  wire [2:0] v_8737_0;
  wire [2:0] v_8738_0;
  wire [2:0] v_8739_0;
  wire [2:0] v_8740_0;
  wire [2:0] v_8741_0;
  wire [2:0] v_8742_0;
  wire [2:0] v_8743_0;
  wire [2:0] v_8744_0;
  wire [2:0] v_8745_0;
  wire [2:0] v_8746_0;
  wire [2:0] v_8747_0;
  wire [2:0] v_8748_0;
  wire [2:0] v_8749_0;
  wire [2:0] v_8750_0;
  wire [2:0] v_8751_0;
  wire [2:0] v_8752_0;
  wire [2:0] v_8753_0;
  wire [2:0] v_8754_0;
  wire [2:0] v_8755_0;
  wire [2:0] v_8756_0;
  wire [2:0] v_8757_0;
  wire [2:0] v_8758_0;
  wire [2:0] v_8759_0;
  wire [2:0] v_8760_0;
  wire [2:0] v_8761_0;
  wire [2:0] v_8762_0;
  wire [2:0] v_8763_0;
  wire [2:0] v_8764_0;
  wire [2:0] v_8765_0;
  wire [2:0] v_8766_0;
  wire [2:0] v_8767_0;
  wire [2:0] v_8768_0;
  wire [2:0] v_8769_0;
  wire [2:0] v_8770_0;
  wire [2:0] v_8771_0;
  wire [2:0] v_8772_0;
  wire [2:0] v_8773_0;
  wire [2:0] v_8774_0;
  wire [2:0] v_8775_0;
  wire [2:0] v_8776_0;
  wire [2:0] v_8777_0;
  wire [2:0] v_8778_0;
  wire [2:0] v_8779_0;
  wire [2:0] v_8780_0;
  wire [2:0] v_8781_0;
  wire [2:0] v_8782_0;
  wire [2:0] v_8783_0;
  wire [2:0] v_8784_0;
  wire [2:0] v_8785_0;
  wire [2:0] v_8786_0;
  wire [2:0] v_8787_0;
  wire [2:0] v_8788_0;
  wire [2:0] v_8789_0;
  wire [2:0] v_8790_0;
  wire [2:0] v_8791_0;
  wire [2:0] v_8792_0;
  wire [2:0] v_8793_0;
  wire [2:0] v_8794_0;
  wire [2:0] v_8795_0;
  wire [2:0] v_8796_0;
  wire [2:0] v_8797_0;
  wire [2:0] v_8798_0;
  wire [2:0] v_8799_0;
  wire [2:0] v_8800_0;
  wire [2:0] v_8801_0;
  wire [2:0] v_8802_0;
  wire [2:0] v_8803_0;
  wire [2:0] v_8804_0;
  wire [2:0] v_8805_0;
  wire [2:0] v_8806_0;
  wire [2:0] v_8807_0;
  wire [2:0] v_8808_0;
  wire [2:0] v_8809_0;
  wire [2:0] v_8810_0;
  wire [2:0] v_8811_0;
  wire [2:0] v_8812_0;
  wire [2:0] v_8813_0;
  wire [2:0] v_8814_0;
  wire [2:0] v_8815_0;
  wire [2:0] v_8816_0;
  wire [2:0] v_8817_0;
  wire [2:0] v_8818_0;
  wire [2:0] v_8819_0;
  wire [2:0] v_8820_0;
  wire [2:0] v_8821_0;
  wire [2:0] v_8822_0;
  wire [2:0] v_8823_0;
  wire [2:0] v_8824_0;
  wire [2:0] v_8825_0;
  wire [2:0] v_8826_0;
  wire [2:0] v_8827_0;
  wire [2:0] v_8828_0;
  wire [2:0] v_8829_0;
  wire [2:0] v_8830_0;
  wire [2:0] v_8831_0;
  wire [2:0] v_8832_0;
  wire [2:0] v_8833_0;
  wire [2:0] v_8834_0;
  wire [2:0] v_8835_0;
  wire [2:0] v_8836_0;
  wire [2:0] v_8837_0;
  wire [2:0] v_8838_0;
  wire [2:0] v_8839_0;
  wire [2:0] v_8840_0;
  wire [2:0] v_8841_0;
  wire [2:0] v_8842_0;
  wire [2:0] v_8843_0;
  wire [2:0] v_8844_0;
  wire [2:0] v_8845_0;
  wire [2:0] v_8846_0;
  wire [2:0] v_8847_0;
  wire [2:0] v_8848_0;
  wire [2:0] v_8849_0;
  wire [2:0] v_8850_0;
  wire [2:0] v_8851_0;
  wire [2:0] v_8852_0;
  wire [2:0] v_8853_0;
  wire [2:0] v_8854_0;
  wire [2:0] v_8855_0;
  wire [2:0] v_8856_0;
  wire [2:0] v_8857_0;
  wire [2:0] v_8858_0;
  wire [2:0] v_8859_0;
  wire [2:0] v_8860_0;
  wire [2:0] v_8861_0;
  wire [2:0] v_8862_0;
  wire [2:0] v_8863_0;
  wire [2:0] v_8864_0;
  wire [2:0] v_8865_0;
  wire [2:0] v_8866_0;
  wire [2:0] v_8867_0;
  wire [2:0] v_8868_0;
  wire [2:0] v_8869_0;
  wire [2:0] v_8870_0;
  wire [2:0] v_8871_0;
  wire [2:0] v_8872_0;
  wire [2:0] v_8873_0;
  wire [2:0] v_8874_0;
  wire [2:0] v_8875_0;
  wire [2:0] v_8876_0;
  wire [2:0] v_8877_0;
  wire [2:0] v_8878_0;
  wire [2:0] v_8879_0;
  wire [2:0] v_8880_0;
  wire [2:0] v_8881_0;
  wire [2:0] v_8882_0;
  wire [2:0] v_8883_0;
  wire [2:0] v_8884_0;
  wire [2:0] v_8885_0;
  wire [2:0] v_8886_0;
  wire [2:0] v_8887_0;
  wire [2:0] v_8888_0;
  wire [2:0] v_8889_0;
  wire [2:0] v_8890_0;
  wire [2:0] v_8891_0;
  wire [2:0] v_8892_0;
  wire [2:0] v_8893_0;
  wire [2:0] v_8894_0;
  wire [2:0] v_8895_0;
  wire [2:0] v_8896_0;
  wire [2:0] v_8897_0;
  wire [2:0] v_8898_0;
  wire [2:0] v_8899_0;
  wire [2:0] v_8900_0;
  wire [2:0] v_8901_0;
  wire [2:0] v_8902_0;
  wire [2:0] v_8903_0;
  wire [2:0] v_8904_0;
  wire [2:0] v_8905_0;
  wire [2:0] v_8906_0;
  wire [2:0] v_8907_0;
  wire [2:0] v_8908_0;
  wire [2:0] v_8909_0;
  wire [2:0] v_8910_0;
  wire [2:0] v_8911_0;
  wire [2:0] v_8912_0;
  wire [2:0] v_8913_0;
  wire [2:0] v_8914_0;
  wire [2:0] v_8915_0;
  wire [2:0] v_8916_0;
  wire [2:0] v_8917_0;
  wire [2:0] v_8918_0;
  wire [2:0] v_8919_0;
  wire [2:0] v_8920_0;
  wire [2:0] v_8921_0;
  wire [2:0] v_8922_0;
  wire [2:0] v_8923_0;
  wire [2:0] v_8924_0;
  wire [2:0] v_8925_0;
  wire [2:0] v_8926_0;
  wire [2:0] v_8927_0;
  wire [2:0] v_8928_0;
  wire [2:0] v_8929_0;
  wire [2:0] v_8930_0;
  wire [2:0] v_8931_0;
  wire [2:0] v_8932_0;
  wire [2:0] v_8933_0;
  wire [2:0] v_8934_0;
  wire [2:0] v_8935_0;
  wire [2:0] v_8936_0;
  wire [2:0] v_8937_0;
  wire [2:0] v_8938_0;
  wire [2:0] v_8939_0;
  wire [2:0] v_8940_0;
  wire [2:0] v_8941_0;
  wire [2:0] v_8942_0;
  wire [2:0] v_8943_0;
  wire [2:0] v_8944_0;
  wire [2:0] v_8945_0;
  wire [2:0] v_8946_0;
  wire [2:0] v_8947_0;
  wire [2:0] v_8948_0;
  wire [2:0] v_8949_0;
  wire [2:0] v_8950_0;
  wire [2:0] v_8951_0;
  wire [2:0] v_8952_0;
  wire [2:0] v_8953_0;
  wire [2:0] v_8954_0;
  wire [2:0] v_8955_0;
  wire [2:0] v_8956_0;
  wire [2:0] v_8957_0;
  wire [2:0] v_8958_0;
  wire [2:0] v_8959_0;
  wire [2:0] v_8960_0;
  wire [2:0] v_8961_0;
  wire [2:0] v_8962_0;
  wire [2:0] v_8963_0;
  wire [2:0] v_8964_0;
  wire [2:0] v_8965_0;
  wire [2:0] v_8966_0;
  wire [2:0] v_8967_0;
  wire [2:0] v_8968_0;
  wire [2:0] v_8969_0;
  wire [2:0] v_8970_0;
  wire [2:0] v_8971_0;
  wire [2:0] v_8972_0;
  wire [2:0] v_8973_0;
  wire [2:0] v_8974_0;
  wire [2:0] v_8975_0;
  wire [2:0] v_8976_0;
  wire [2:0] v_8977_0;
  wire [2:0] v_8978_0;
  wire [2:0] v_8979_0;
  wire [2:0] v_8980_0;
  wire [2:0] v_8981_0;
  wire [2:0] v_8982_0;
  wire [2:0] v_8983_0;
  wire [2:0] v_8984_0;
  wire [2:0] v_8985_0;
  wire [2:0] v_8986_0;
  wire [2:0] v_8987_0;
  wire [2:0] v_8988_0;
  wire [2:0] v_8989_0;
  wire [2:0] v_8990_0;
  wire [2:0] v_8991_0;
  wire [2:0] v_8992_0;
  wire [2:0] v_8993_0;
  wire [2:0] v_8994_0;
  wire [2:0] v_8995_0;
  wire [2:0] v_8996_0;
  wire [2:0] v_8997_0;
  wire [2:0] v_8998_0;
  wire [2:0] v_8999_0;
  wire [2:0] v_9000_0;
  wire [2:0] v_9001_0;
  wire [2:0] v_9002_0;
  wire [2:0] v_9003_0;
  wire [2:0] v_9004_0;
  wire [2:0] v_9005_0;
  wire [2:0] v_9006_0;
  wire [2:0] v_9007_0;
  wire [2:0] v_9008_0;
  wire [2:0] v_9009_0;
  wire [2:0] v_9010_0;
  wire [2:0] v_9011_0;
  wire [2:0] v_9012_0;
  wire [2:0] v_9013_0;
  wire [2:0] v_9014_0;
  wire [2:0] v_9015_0;
  wire [2:0] v_9016_0;
  wire [2:0] v_9017_0;
  wire [2:0] v_9018_0;
  wire [2:0] v_9019_0;
  wire [2:0] v_9020_0;
  wire [2:0] v_9021_0;
  wire [2:0] v_9022_0;
  wire [2:0] v_9023_0;
  wire [2:0] v_9024_0;
  wire [2:0] v_9025_0;
  wire [2:0] v_9026_0;
  wire [2:0] v_9027_0;
  wire [2:0] v_9028_0;
  wire [2:0] v_9029_0;
  wire [2:0] v_9030_0;
  wire [2:0] v_9031_0;
  wire [2:0] v_9032_0;
  wire [2:0] v_9033_0;
  wire [2:0] v_9034_0;
  wire [2:0] v_9035_0;
  wire [2:0] v_9036_0;
  wire [2:0] v_9037_0;
  wire [2:0] v_9038_0;
  wire [2:0] v_9039_0;
  wire [2:0] v_9040_0;
  wire [2:0] v_9041_0;
  wire [2:0] v_9042_0;
  wire [2:0] v_9043_0;
  wire [2:0] v_9044_0;
  wire [2:0] v_9045_0;
  wire [2:0] v_9046_0;
  wire [2:0] v_9047_0;
  wire [2:0] v_9048_0;
  wire [2:0] v_9049_0;
  wire [2:0] v_9050_0;
  wire [2:0] v_9051_0;
  wire [2:0] v_9052_0;
  wire [2:0] v_9053_0;
  wire [2:0] v_9054_0;
  wire [2:0] v_9055_0;
  wire [2:0] v_9056_0;
  wire [2:0] v_9057_0;
  wire [2:0] v_9058_0;
  wire [2:0] v_9059_0;
  wire [2:0] v_9060_0;
  wire [2:0] v_9061_0;
  wire [2:0] v_9062_0;
  wire [2:0] v_9063_0;
  wire [2:0] v_9064_0;
  wire [2:0] v_9065_0;
  wire [2:0] v_9066_0;
  wire [2:0] v_9067_0;
  wire [2:0] v_9068_0;
  wire [2:0] v_9069_0;
  wire [2:0] v_9070_0;
  wire [2:0] v_9071_0;
  wire [2:0] v_9072_0;
  wire [2:0] v_9073_0;
  wire [2:0] v_9074_0;
  wire [2:0] v_9075_0;
  wire [2:0] v_9076_0;
  wire [2:0] v_9077_0;
  wire [2:0] v_9078_0;
  wire [2:0] v_9079_0;
  wire [2:0] v_9080_0;
  wire [2:0] v_9081_0;
  wire [2:0] v_9082_0;
  wire [2:0] v_9083_0;
  wire [2:0] v_9084_0;
  wire [2:0] v_9085_0;
  wire [2:0] v_9086_0;
  wire [2:0] v_9087_0;
  wire [2:0] v_9088_0;
  wire [2:0] v_9089_0;
  wire [2:0] v_9090_0;
  wire [2:0] v_9091_0;
  wire [2:0] v_9092_0;
  wire [2:0] v_9093_0;
  wire [2:0] v_9094_0;
  wire [2:0] v_9095_0;
  wire [2:0] v_9096_0;
  wire [2:0] v_9097_0;
  wire [2:0] v_9098_0;
  wire [2:0] v_9099_0;
  wire [2:0] v_9100_0;
  wire [2:0] v_9101_0;
  wire [2:0] v_9102_0;
  wire [2:0] v_9103_0;
  wire [2:0] v_9104_0;
  wire [2:0] v_9105_0;
  wire [2:0] v_9106_0;
  wire [2:0] v_9107_0;
  wire [2:0] v_9108_0;
  wire [2:0] v_9109_0;
  wire [2:0] v_9110_0;
  wire [2:0] v_9111_0;
  wire [2:0] v_9112_0;
  wire [2:0] v_9113_0;
  wire [2:0] v_9114_0;
  wire [2:0] v_9115_0;
  wire [2:0] v_9116_0;
  wire [2:0] v_9117_0;
  wire [2:0] v_9118_0;
  wire [2:0] v_9119_0;
  wire [2:0] v_9120_0;
  wire [2:0] v_9121_0;
  wire [2:0] v_9122_0;
  wire [2:0] v_9123_0;
  wire [2:0] v_9124_0;
  wire [2:0] v_9125_0;
  wire [2:0] v_9126_0;
  wire [2:0] v_9127_0;
  wire [2:0] v_9128_0;
  wire [2:0] v_9129_0;
  wire [2:0] v_9130_0;
  wire [2:0] v_9131_0;
  wire [2:0] v_9132_0;
  wire [2:0] v_9133_0;
  wire [2:0] v_9134_0;
  wire [2:0] v_9135_0;
  wire [2:0] v_9136_0;
  wire [2:0] v_9137_0;
  wire [2:0] v_9138_0;
  wire [2:0] v_9139_0;
  wire [2:0] v_9140_0;
  wire [2:0] v_9141_0;
  wire [2:0] v_9142_0;
  wire [2:0] v_9143_0;
  wire [2:0] v_9144_0;
  wire [2:0] v_9145_0;
  wire [2:0] v_9146_0;
  wire [2:0] v_9147_0;
  wire [2:0] v_9148_0;
  wire [2:0] v_9149_0;
  wire [2:0] v_9150_0;
  wire [2:0] v_9151_0;
  wire [2:0] v_9152_0;
  wire [2:0] v_9153_0;
  wire [2:0] v_9154_0;
  wire [2:0] v_9155_0;
  wire [2:0] v_9156_0;
  wire [2:0] v_9157_0;
  wire [2:0] v_9158_0;
  wire [2:0] v_9159_0;
  wire [2:0] v_9160_0;
  wire [2:0] v_9161_0;
  wire [2:0] v_9162_0;
  wire [2:0] v_9163_0;
  wire [2:0] v_9164_0;
  wire [2:0] v_9165_0;
  wire [2:0] v_9166_0;
  wire [2:0] v_9167_0;
  wire [2:0] v_9168_0;
  wire [2:0] v_9169_0;
  wire [2:0] v_9170_0;
  wire [2:0] v_9171_0;
  wire [2:0] v_9172_0;
  wire [2:0] v_9173_0;
  wire [2:0] v_9174_0;
  wire [2:0] v_9175_0;
  wire [2:0] v_9176_0;
  wire [2:0] v_9177_0;
  wire [2:0] v_9178_0;
  wire [2:0] v_9179_0;
  wire [2:0] v_9180_0;
  wire [2:0] v_9181_0;
  wire [2:0] v_9182_0;
  wire [2:0] v_9183_0;
  wire [2:0] v_9184_0;
  wire [2:0] v_9185_0;
  wire [2:0] v_9186_0;
  wire [2:0] v_9187_0;
  wire [2:0] v_9188_0;
  wire [2:0] v_9189_0;
  wire [2:0] v_9190_0;
  wire [2:0] v_9191_0;
  wire [2:0] v_9192_0;
  wire [2:0] v_9193_0;
  wire [2:0] v_9194_0;
  wire [2:0] v_9195_0;
  wire [2:0] v_9196_0;
  wire [2:0] v_9197_0;
  wire [2:0] v_9198_0;
  wire [2:0] v_9199_0;
  wire [2:0] v_9200_0;
  wire [2:0] v_9201_0;
  wire [2:0] v_9202_0;
  wire [2:0] v_9203_0;
  wire [2:0] v_9204_0;
  wire [2:0] v_9205_0;
  wire [2:0] v_9206_0;
  wire [2:0] v_9207_0;
  wire [2:0] v_9208_0;
  wire [2:0] v_9209_0;
  wire [2:0] v_9210_0;
  wire [2:0] v_9211_0;
  wire [2:0] v_9212_0;
  wire [2:0] v_9213_0;
  wire [2:0] v_9214_0;
  wire [2:0] v_9215_0;
  wire [2:0] v_9216_0;
  wire [2:0] v_9217_0;
  wire [2:0] v_9218_0;
  wire [2:0] v_9219_0;
  wire [2:0] v_9220_0;
  wire [2:0] v_9221_0;
  wire [2:0] v_9222_0;
  wire [2:0] v_9223_0;
  wire [2:0] v_9224_0;
  wire [2:0] v_9225_0;
  wire [2:0] v_9226_0;
  wire [2:0] v_9227_0;
  wire [2:0] v_9228_0;
  wire [2:0] v_9229_0;
  wire [2:0] v_9230_0;
  wire [2:0] v_9231_0;
  wire [2:0] v_9232_0;
  wire [2:0] v_9233_0;
  wire [2:0] v_9234_0;
  wire [2:0] v_9235_0;
  wire [2:0] v_9236_0;
  wire [2:0] v_9237_0;
  wire [2:0] v_9238_0;
  wire [2:0] v_9239_0;
  wire [2:0] v_9240_0;
  wire [2:0] v_9241_0;
  wire [2:0] v_9242_0;
  wire [2:0] v_9243_0;
  wire [2:0] v_9244_0;
  wire [2:0] v_9245_0;
  wire [2:0] v_9246_0;
  wire [2:0] v_9247_0;
  wire [2:0] v_9248_0;
  wire [2:0] v_9249_0;
  wire [2:0] v_9250_0;
  wire [2:0] v_9251_0;
  wire [2:0] v_9252_0;
  wire [2:0] v_9253_0;
  wire [2:0] v_9254_0;
  wire [2:0] v_9255_0;
  wire [2:0] v_9256_0;
  wire [2:0] v_9257_0;
  wire [2:0] v_9258_0;
  wire [2:0] v_9259_0;
  wire [2:0] v_9260_0;
  wire [2:0] v_9261_0;
  wire [2:0] v_9262_0;
  wire [2:0] v_9263_0;
  wire [2:0] v_9264_0;
  wire [2:0] v_9265_0;
  wire [2:0] v_9266_0;
  wire [2:0] v_9267_0;
  wire [2:0] v_9268_0;
  wire [2:0] v_9269_0;
  wire [2:0] v_9270_0;
  wire [2:0] v_9271_0;
  wire [2:0] v_9272_0;
  wire [2:0] v_9273_0;
  wire [2:0] v_9274_0;
  wire [2:0] v_9275_0;
  wire [2:0] v_9276_0;
  wire [2:0] v_9277_0;
  wire [2:0] v_9278_0;
  wire [2:0] v_9279_0;
  wire [2:0] v_9280_0;
  wire [2:0] v_9281_0;
  wire [2:0] v_9282_0;
  wire [2:0] v_9283_0;
  wire [2:0] v_9284_0;
  wire [2:0] v_9285_0;
  wire [2:0] v_9286_0;
  wire [2:0] v_9287_0;
  wire [2:0] v_9288_0;
  wire [2:0] v_9289_0;
  wire [2:0] v_9290_0;
  wire [2:0] v_9291_0;
  wire [2:0] v_9292_0;
  wire [2:0] v_9293_0;
  wire [2:0] v_9294_0;
  wire [2:0] v_9295_0;
  wire [2:0] v_9296_0;
  wire [2:0] v_9297_0;
  wire [2:0] v_9298_0;
  wire [2:0] v_9299_0;
  wire [2:0] v_9300_0;
  wire [2:0] v_9301_0;
  wire [2:0] v_9302_0;
  wire [2:0] v_9303_0;
  wire [2:0] v_9304_0;
  wire [2:0] v_9305_0;
  wire [2:0] v_9306_0;
  wire [2:0] v_9307_0;
  wire [2:0] v_9308_0;
  wire [2:0] v_9309_0;
  wire [2:0] v_9310_0;
  wire [2:0] v_9311_0;
  wire [2:0] v_9312_0;
  wire [2:0] v_9313_0;
  wire [2:0] v_9314_0;
  wire [2:0] v_9315_0;
  wire [2:0] v_9316_0;
  wire [2:0] v_9317_0;
  wire [2:0] v_9318_0;
  wire [2:0] v_9319_0;
  wire [2:0] v_9320_0;
  wire [2:0] v_9321_0;
  wire [2:0] v_9322_0;
  wire [2:0] v_9323_0;
  wire [2:0] v_9324_0;
  wire [2:0] v_9325_0;
  wire [2:0] v_9326_0;
  wire [2:0] v_9327_0;
  wire [2:0] v_9328_0;
  wire [2:0] v_9329_0;
  wire [2:0] v_9330_0;
  wire [2:0] v_9331_0;
  wire [2:0] v_9332_0;
  wire [2:0] v_9333_0;
  wire [2:0] v_9334_0;
  wire [2:0] v_9335_0;
  wire [2:0] v_9336_0;
  wire [2:0] v_9337_0;
  wire [2:0] v_9338_0;
  wire [2:0] v_9339_0;
  wire [2:0] v_9340_0;
  wire [2:0] v_9341_0;
  wire [2:0] v_9342_0;
  wire [2:0] v_9343_0;
  wire [2:0] v_9344_0;
  wire [2:0] v_9345_0;
  wire [2:0] v_9346_0;
  wire [2:0] v_9347_0;
  wire [2:0] v_9348_0;
  wire [2:0] v_9349_0;
  wire [2:0] v_9350_0;
  wire [2:0] v_9351_0;
  wire [2:0] v_9352_0;
  wire [2:0] v_9353_0;
  wire [2:0] v_9354_0;
  wire [2:0] v_9355_0;
  wire [2:0] v_9356_0;
  wire [2:0] v_9357_0;
  wire [2:0] v_9358_0;
  wire [2:0] v_9359_0;
  wire [2:0] v_9360_0;
  wire [2:0] v_9361_0;
  wire [2:0] v_9362_0;
  wire [2:0] v_9363_0;
  wire [2:0] v_9364_0;
  wire [2:0] v_9365_0;
  wire [2:0] v_9366_0;
  wire [2:0] v_9367_0;
  wire [2:0] v_9368_0;
  wire [2:0] v_9369_0;
  wire [2:0] v_9370_0;
  wire [2:0] v_9371_0;
  wire [2:0] v_9372_0;
  wire [2:0] v_9373_0;
  wire [2:0] v_9374_0;
  wire [2:0] v_9375_0;
  wire [2:0] v_9376_0;
  wire [2:0] v_9377_0;
  wire [2:0] v_9378_0;
  wire [2:0] v_9379_0;
  wire [2:0] v_9380_0;
  wire [2:0] v_9381_0;
  wire [2:0] v_9382_0;
  wire [2:0] v_9383_0;
  wire [2:0] v_9384_0;
  wire [2:0] v_9385_0;
  wire [2:0] v_9386_0;
  wire [2:0] v_9387_0;
  wire [2:0] v_9388_0;
  wire [2:0] v_9389_0;
  wire [2:0] v_9390_0;
  wire [2:0] v_9391_0;
  wire [2:0] v_9392_0;
  wire [2:0] v_9393_0;
  wire [2:0] v_9394_0;
  wire [2:0] v_9395_0;
  wire [2:0] v_9396_0;
  wire [2:0] v_9397_0;
  wire [2:0] v_9398_0;
  wire [2:0] v_9399_0;
  wire [2:0] v_9400_0;
  wire [2:0] v_9401_0;
  wire [2:0] v_9402_0;
  wire [2:0] v_9403_0;
  wire [2:0] v_9404_0;
  wire [2:0] v_9405_0;
  wire [2:0] v_9406_0;
  wire [2:0] v_9407_0;
  wire [2:0] v_9408_0;
  wire [2:0] v_9409_0;
  wire [2:0] v_9410_0;
  wire [2:0] v_9411_0;
  wire [2:0] v_9412_0;
  wire [2:0] v_9413_0;
  wire [2:0] v_9414_0;
  wire [2:0] v_9415_0;
  wire [2:0] v_9416_0;
  wire [2:0] v_9417_0;
  wire [2:0] v_9418_0;
  wire [2:0] v_9419_0;
  wire [2:0] v_9420_0;
  wire [2:0] v_9421_0;
  wire [2:0] v_9422_0;
  wire [2:0] v_9423_0;
  wire [2:0] v_9424_0;
  wire [2:0] v_9425_0;
  wire [2:0] v_9426_0;
  wire [2:0] v_9427_0;
  wire [2:0] v_9428_0;
  wire [2:0] v_9429_0;
  wire [2:0] v_9430_0;
  wire [2:0] v_9431_0;
  wire [2:0] v_9432_0;
  wire [2:0] v_9433_0;
  wire [2:0] v_9434_0;
  wire [2:0] v_9435_0;
  wire [2:0] v_9436_0;
  wire [2:0] v_9437_0;
  wire [2:0] v_9438_0;
  wire [2:0] v_9439_0;
  wire [2:0] v_9440_0;
  wire [2:0] v_9441_0;
  wire [2:0] v_9442_0;
  wire [2:0] v_9443_0;
  wire [2:0] v_9444_0;
  wire [2:0] v_9445_0;
  wire [2:0] v_9446_0;
  wire [2:0] v_9447_0;
  wire [2:0] v_9448_0;
  wire [2:0] v_9449_0;
  wire [2:0] v_9450_0;
  wire [2:0] v_9451_0;
  wire [2:0] v_9452_0;
  wire [2:0] v_9453_0;
  wire [2:0] v_9454_0;
  wire [2:0] v_9455_0;
  wire [2:0] v_9456_0;
  wire [2:0] v_9457_0;
  wire [2:0] v_9458_0;
  wire [2:0] v_9459_0;
  wire [2:0] v_9460_0;
  wire [2:0] v_9461_0;
  wire [2:0] v_9462_0;
  wire [2:0] v_9463_0;
  wire [2:0] v_9464_0;
  wire [2:0] v_9465_0;
  wire [2:0] v_9466_0;
  wire [2:0] v_9467_0;
  wire [2:0] v_9468_0;
  wire [2:0] v_9469_0;
  wire [2:0] v_9470_0;
  wire [2:0] v_9471_0;
  wire [2:0] v_9472_0;
  wire [2:0] v_9473_0;
  wire [2:0] v_9474_0;
  wire [2:0] v_9475_0;
  wire [2:0] v_9476_0;
  wire [2:0] v_9477_0;
  wire [2:0] v_9478_0;
  wire [2:0] v_9479_0;
  wire [2:0] v_9480_0;
  wire [2:0] v_9481_0;
  wire [2:0] v_9482_0;
  wire [2:0] v_9483_0;
  wire [2:0] v_9484_0;
  wire [2:0] v_9485_0;
  wire [2:0] v_9486_0;
  wire [2:0] v_9487_0;
  wire [2:0] v_9488_0;
  wire [2:0] v_9489_0;
  wire [2:0] v_9490_0;
  wire [2:0] v_9491_0;
  wire [2:0] v_9492_0;
  wire [2:0] v_9493_0;
  wire [2:0] v_9494_0;
  wire [2:0] v_9495_0;
  wire [2:0] v_9496_0;
  wire [2:0] v_9497_0;
  wire [2:0] v_9498_0;
  wire [2:0] v_9499_0;
  wire [2:0] v_9500_0;
  wire [2:0] v_9501_0;
  wire [2:0] v_9502_0;
  wire [2:0] v_9503_0;
  wire [2:0] v_9504_0;
  wire [2:0] v_9505_0;
  wire [2:0] v_9506_0;
  wire [2:0] v_9507_0;
  wire [2:0] v_9508_0;
  wire [2:0] v_9509_0;
  wire [2:0] v_9510_0;
  wire [2:0] v_9511_0;
  wire [2:0] v_9512_0;
  wire [2:0] v_9513_0;
  wire [2:0] v_9514_0;
  wire [2:0] v_9515_0;
  wire [2:0] v_9516_0;
  wire [2:0] v_9517_0;
  wire [2:0] v_9518_0;
  wire [2:0] v_9519_0;
  wire [2:0] v_9520_0;
  wire [2:0] v_9521_0;
  wire [2:0] v_9522_0;
  wire [2:0] v_9523_0;
  wire [2:0] v_9524_0;
  wire [2:0] v_9525_0;
  wire [2:0] v_9526_0;
  wire [2:0] v_9527_0;
  wire [2:0] v_9528_0;
  wire [2:0] v_9529_0;
  wire [2:0] v_9530_0;
  wire [2:0] v_9531_0;
  wire [2:0] v_9532_0;
  wire [2:0] v_9533_0;
  wire [2:0] v_9534_0;
  wire [2:0] v_9535_0;
  wire [2:0] v_9536_0;
  wire [2:0] v_9537_0;
  wire [2:0] v_9538_0;
  wire [2:0] v_9539_0;
  wire [2:0] v_9540_0;
  wire [2:0] v_9541_0;
  wire [2:0] v_9542_0;
  wire [2:0] v_9543_0;
  wire [2:0] v_9544_0;
  wire [2:0] v_9545_0;
  wire [2:0] v_9546_0;
  wire [2:0] v_9547_0;
  wire [2:0] v_9548_0;
  wire [2:0] v_9549_0;
  wire [2:0] v_9550_0;
  wire [2:0] v_9551_0;
  wire [2:0] v_9552_0;
  wire [2:0] v_9553_0;
  wire [2:0] v_9554_0;
  wire [2:0] v_9555_0;
  wire [2:0] v_9556_0;
  wire [2:0] v_9557_0;
  wire [2:0] v_9558_0;
  wire [2:0] v_9559_0;
  wire [2:0] v_9560_0;
  wire [2:0] v_9561_0;
  wire [2:0] v_9562_0;
  wire [2:0] v_9563_0;
  wire [2:0] v_9564_0;
  wire [2:0] v_9565_0;
  wire [2:0] v_9566_0;
  wire [2:0] v_9567_0;
  wire [2:0] v_9568_0;
  wire [2:0] v_9569_0;
  wire [2:0] v_9570_0;
  wire [2:0] v_9571_0;
  wire [2:0] v_9572_0;
  wire [2:0] v_9573_0;
  wire [2:0] v_9574_0;
  wire [2:0] v_9575_0;
  wire [2:0] v_9576_0;
  wire [2:0] v_9577_0;
  wire [2:0] v_9578_0;
  wire [2:0] v_9579_0;
  wire [2:0] v_9580_0;
  wire [2:0] v_9581_0;
  wire [2:0] v_9582_0;
  wire [2:0] v_9583_0;
  wire [2:0] v_9584_0;
  wire [2:0] v_9585_0;
  wire [2:0] v_9586_0;
  wire [2:0] v_9587_0;
  wire [2:0] v_9588_0;
  wire [2:0] v_9589_0;
  wire [2:0] v_9590_0;
  wire [2:0] v_9591_0;
  wire [2:0] v_9592_0;
  wire [2:0] v_9593_0;
  wire [2:0] v_9594_0;
  wire [2:0] v_9595_0;
  wire [2:0] v_9596_0;
  wire [2:0] v_9597_0;
  wire [2:0] v_9598_0;
  wire [2:0] v_9599_0;
  wire [2:0] v_9600_0;
  wire [2:0] v_9601_0;
  wire [2:0] v_9602_0;
  wire [2:0] v_9603_0;
  wire [2:0] v_9604_0;
  wire [2:0] v_9605_0;
  wire [2:0] v_9606_0;
  wire [2:0] v_9607_0;
  wire [2:0] v_9608_0;
  wire [2:0] v_9609_0;
  wire [2:0] v_9610_0;
  wire [2:0] v_9611_0;
  wire [2:0] v_9612_0;
  wire [2:0] v_9613_0;
  wire [2:0] v_9614_0;
  wire [2:0] v_9615_0;
  wire [2:0] v_9616_0;
  wire [2:0] v_9617_0;
  wire [2:0] v_9618_0;
  wire [2:0] v_9619_0;
  wire [2:0] v_9620_0;
  wire [2:0] v_9621_0;
  wire [2:0] v_9622_0;
  wire [2:0] v_9623_0;
  wire [2:0] v_9624_0;
  wire [2:0] v_9625_0;
  wire [2:0] v_9626_0;
  wire [2:0] v_9627_0;
  wire [2:0] v_9628_0;
  wire [2:0] v_9629_0;
  wire [2:0] v_9630_0;
  wire [2:0] v_9631_0;
  wire [2:0] v_9632_0;
  wire [2:0] v_9633_0;
  wire [2:0] v_9634_0;
  wire [2:0] v_9635_0;
  wire [2:0] v_9636_0;
  wire [2:0] v_9637_0;
  wire [2:0] v_9638_0;
  wire [2:0] v_9639_0;
  wire [2:0] v_9640_0;
  wire [2:0] v_9641_0;
  wire [2:0] v_9642_0;
  wire [2:0] v_9643_0;
  wire [2:0] v_9644_0;
  wire [2:0] v_9645_0;
  wire [2:0] v_9646_0;
  wire [2:0] v_9647_0;
  wire [2:0] v_9648_0;
  wire [2:0] v_9649_0;
  wire [2:0] v_9650_0;
  wire [2:0] v_9651_0;
  wire [2:0] v_9652_0;
  wire [2:0] v_9653_0;
  wire [2:0] v_9654_0;
  wire [2:0] v_9655_0;
  wire [2:0] v_9656_0;
  wire [2:0] v_9657_0;
  wire [2:0] v_9658_0;
  wire [2:0] v_9659_0;
  wire [2:0] v_9660_0;
  wire [2:0] v_9661_0;
  wire [2:0] v_9662_0;
  wire [2:0] v_9663_0;
  wire [2:0] v_9664_0;
  wire [2:0] v_9665_0;
  wire [2:0] v_9666_0;
  wire [2:0] v_9667_0;
  wire [2:0] v_9668_0;
  wire [2:0] v_9669_0;
  wire [2:0] v_9670_0;
  wire [2:0] v_9671_0;
  wire [2:0] v_9672_0;
  wire [2:0] v_9673_0;
  wire [2:0] v_9674_0;
  wire [2:0] v_9675_0;
  wire [2:0] v_9676_0;
  wire [2:0] v_9677_0;
  wire [2:0] v_9678_0;
  wire [2:0] v_9679_0;
  wire [2:0] v_9680_0;
  wire [2:0] v_9681_0;
  wire [2:0] v_9682_0;
  wire [2:0] v_9683_0;
  wire [2:0] v_9684_0;
  wire [2:0] v_9685_0;
  wire [2:0] v_9686_0;
  wire [2:0] v_9687_0;
  wire [2:0] v_9688_0;
  wire [2:0] v_9689_0;
  wire [2:0] v_9690_0;
  wire [2:0] v_9691_0;
  wire [2:0] v_9692_0;
  wire [2:0] v_9693_0;
  wire [2:0] v_9694_0;
  wire [2:0] v_9695_0;
  wire [2:0] v_9696_0;
  wire [2:0] v_9697_0;
  wire [2:0] v_9698_0;
  wire [2:0] v_9699_0;
  wire [2:0] v_9700_0;
  wire [2:0] v_9701_0;
  wire [2:0] v_9702_0;
  wire [2:0] v_9703_0;
  wire [2:0] v_9704_0;
  wire [2:0] v_9705_0;
  wire [2:0] v_9706_0;
  wire [2:0] v_9707_0;
  wire [2:0] v_9708_0;
  wire [2:0] v_9709_0;
  wire [2:0] v_9710_0;
  wire [2:0] v_9711_0;
  wire [2:0] v_9712_0;
  wire [2:0] v_9713_0;
  wire [2:0] v_9714_0;
  wire [2:0] v_9715_0;
  wire [2:0] v_9716_0;
  wire [2:0] v_9717_0;
  wire [2:0] v_9718_0;
  wire [2:0] v_9719_0;
  wire [2:0] v_9720_0;
  wire [2:0] v_9721_0;
  wire [2:0] v_9722_0;
  wire [2:0] v_9723_0;
  wire [2:0] v_9724_0;
  wire [2:0] v_9725_0;
  wire [2:0] v_9726_0;
  wire [2:0] v_9727_0;
  wire [2:0] v_9728_0;
  wire [2:0] v_9729_0;
  wire [2:0] v_9730_0;
  wire [2:0] v_9731_0;
  wire [2:0] v_9732_0;
  wire [2:0] v_9733_0;
  wire [2:0] v_9734_0;
  wire [2:0] v_9735_0;
  wire [2:0] v_9736_0;
  wire [2:0] v_9737_0;
  wire [2:0] v_9738_0;
  wire [2:0] v_9739_0;
  wire [2:0] v_9740_0;
  wire [2:0] v_9741_0;
  wire [2:0] v_9742_0;
  wire [2:0] v_9743_0;
  wire [2:0] v_9744_0;
  wire [2:0] v_9745_0;
  wire [2:0] v_9746_0;
  wire [2:0] v_9747_0;
  wire [2:0] v_9748_0;
  wire [2:0] v_9749_0;
  wire [2:0] v_9750_0;
  wire [2:0] v_9751_0;
  wire [2:0] v_9752_0;
  wire [2:0] v_9753_0;
  wire [2:0] v_9754_0;
  wire [2:0] v_9755_0;
  wire [2:0] v_9756_0;
  wire [2:0] v_9757_0;
  wire [2:0] v_9758_0;
  wire [2:0] v_9759_0;
  wire [2:0] v_9760_0;
  wire [2:0] v_9761_0;
  wire [2:0] v_9762_0;
  wire [2:0] v_9763_0;
  wire [2:0] v_9764_0;
  wire [2:0] v_9765_0;
  wire [2:0] v_9766_0;
  wire [2:0] v_9767_0;
  wire [2:0] v_9768_0;
  wire [2:0] v_9769_0;
  wire [2:0] v_9770_0;
  wire [2:0] v_9771_0;
  wire [2:0] v_9772_0;
  wire [2:0] v_9773_0;
  wire [2:0] v_9774_0;
  wire [2:0] v_9775_0;
  wire [2:0] v_9776_0;
  wire [2:0] v_9777_0;
  wire [2:0] v_9778_0;
  wire [2:0] v_9779_0;
  wire [2:0] v_9780_0;
  wire [2:0] v_9781_0;
  wire [2:0] v_9782_0;
  wire [2:0] v_9783_0;
  wire [2:0] v_9784_0;
  wire [2:0] v_9785_0;
  wire [2:0] v_9786_0;
  wire [2:0] v_9787_0;
  wire [2:0] v_9788_0;
  wire [2:0] v_9789_0;
  wire [2:0] v_9790_0;
  wire [2:0] v_9791_0;
  wire [2:0] v_9792_0;
  wire [2:0] v_9793_0;
  wire [2:0] v_9794_0;
  wire [2:0] v_9795_0;
  wire [2:0] v_9796_0;
  wire [2:0] v_9797_0;
  wire [2:0] v_9798_0;
  wire [2:0] v_9799_0;
  wire [2:0] v_9800_0;
  wire [2:0] v_9801_0;
  wire [2:0] v_9802_0;
  wire [2:0] v_9803_0;
  wire [2:0] v_9804_0;
  wire [2:0] v_9805_0;
  wire [2:0] v_9806_0;
  wire [2:0] v_9807_0;
  wire [2:0] v_9808_0;
  wire [2:0] v_9809_0;
  wire [2:0] v_9810_0;
  wire [2:0] v_9811_0;
  wire [2:0] v_9812_0;
  wire [2:0] v_9813_0;
  wire [2:0] v_9814_0;
  wire [2:0] v_9815_0;
  wire [2:0] v_9816_0;
  wire [2:0] v_9817_0;
  wire [2:0] v_9818_0;
  wire [2:0] v_9819_0;
  wire [2:0] v_9820_0;
  wire [2:0] v_9821_0;
  wire [2:0] v_9822_0;
  wire [2:0] v_9823_0;
  wire [2:0] v_9824_0;
  wire [2:0] v_9825_0;
  wire [2:0] v_9826_0;
  wire [2:0] v_9827_0;
  wire [2:0] v_9828_0;
  wire [2:0] v_9829_0;
  wire [2:0] v_9830_0;
  wire [2:0] v_9831_0;
  wire [2:0] v_9832_0;
  wire [2:0] v_9833_0;
  wire [2:0] v_9834_0;
  wire [2:0] v_9835_0;
  wire [2:0] v_9836_0;
  wire [2:0] v_9837_0;
  wire [2:0] v_9838_0;
  wire [2:0] v_9839_0;
  wire [2:0] v_9840_0;
  wire [2:0] v_9841_0;
  wire [2:0] v_9842_0;
  wire [2:0] v_9843_0;
  wire [2:0] v_9844_0;
  wire [2:0] v_9845_0;
  wire [2:0] v_9846_0;
  wire [2:0] v_9847_0;
  wire [2:0] v_9848_0;
  wire [2:0] v_9849_0;
  wire [2:0] v_9850_0;
  wire [2:0] v_9851_0;
  wire [2:0] v_9852_0;
  wire [2:0] v_9853_0;
  wire [2:0] v_9854_0;
  wire [2:0] v_9855_0;
  wire [2:0] v_9856_0;
  wire [2:0] v_9857_0;
  wire [2:0] v_9858_0;
  wire [2:0] v_9859_0;
  wire [2:0] v_9860_0;
  wire [2:0] v_9861_0;
  wire [2:0] v_9862_0;
  wire [2:0] v_9863_0;
  wire [2:0] v_9864_0;
  wire [2:0] v_9865_0;
  wire [2:0] v_9866_0;
  wire [2:0] v_9867_0;
  wire [2:0] v_9868_0;
  wire [2:0] v_9869_0;
  wire [2:0] v_9870_0;
  wire [2:0] v_9871_0;
  wire [2:0] v_9872_0;
  wire [2:0] v_9873_0;
  wire [2:0] v_9874_0;
  wire [2:0] v_9875_0;
  wire [2:0] v_9876_0;
  wire [2:0] v_9877_0;
  wire [2:0] v_9878_0;
  wire [2:0] v_9879_0;
  wire [2:0] v_9880_0;
  wire [2:0] v_9881_0;
  wire [2:0] v_9882_0;
  wire [2:0] v_9883_0;
  wire [2:0] v_9884_0;
  wire [2:0] v_9885_0;
  wire [2:0] v_9886_0;
  wire [2:0] v_9887_0;
  wire [2:0] v_9888_0;
  wire [2:0] v_9889_0;
  wire [2:0] v_9890_0;
  wire [2:0] v_9891_0;
  wire [2:0] v_9892_0;
  wire [2:0] v_9893_0;
  wire [2:0] v_9894_0;
  wire [2:0] v_9895_0;
  wire [2:0] v_9896_0;
  wire [2:0] v_9897_0;
  wire [2:0] v_9898_0;
  wire [2:0] v_9899_0;
  wire [2:0] v_9900_0;
  wire [2:0] v_9901_0;
  wire [2:0] v_9902_0;
  wire [2:0] v_9903_0;
  wire [2:0] v_9904_0;
  wire [2:0] v_9905_0;
  wire [2:0] v_9906_0;
  wire [2:0] v_9907_0;
  wire [2:0] v_9908_0;
  wire [2:0] v_9909_0;
  wire [2:0] v_9910_0;
  wire [2:0] v_9911_0;
  wire [2:0] v_9912_0;
  wire [2:0] v_9913_0;
  wire [2:0] v_9914_0;
  wire [2:0] v_9915_0;
  wire [2:0] v_9916_0;
  wire [2:0] v_9917_0;
  wire [2:0] v_9918_0;
  wire [2:0] v_9919_0;
  wire [2:0] v_9920_0;
  wire [2:0] v_9921_0;
  wire [2:0] v_9922_0;
  wire [2:0] v_9923_0;
  wire [2:0] v_9924_0;
  wire [2:0] v_9925_0;
  wire [2:0] v_9926_0;
  wire [2:0] v_9927_0;
  wire [2:0] v_9928_0;
  wire [2:0] v_9929_0;
  wire [2:0] v_9930_0;
  wire [2:0] v_9931_0;
  wire [2:0] v_9932_0;
  wire [2:0] v_9933_0;
  wire [2:0] v_9934_0;
  wire [2:0] v_9935_0;
  wire [2:0] v_9936_0;
  wire [2:0] v_9937_0;
  wire [2:0] v_9938_0;
  wire [2:0] v_9939_0;
  wire [2:0] v_9940_0;
  wire [2:0] v_9941_0;
  wire [2:0] v_9942_0;
  wire [2:0] v_9943_0;
  wire [2:0] v_9944_0;
  wire [2:0] v_9945_0;
  wire [2:0] v_9946_0;
  wire [2:0] v_9947_0;
  wire [2:0] v_9948_0;
  wire [2:0] v_9949_0;
  wire [2:0] v_9950_0;
  wire [2:0] v_9951_0;
  wire [2:0] v_9952_0;
  wire [2:0] v_9953_0;
  wire [2:0] v_9954_0;
  wire [2:0] v_9955_0;
  wire [2:0] v_9956_0;
  wire [2:0] v_9957_0;
  wire [2:0] v_9958_0;
  wire [2:0] v_9959_0;
  wire [2:0] v_9960_0;
  wire [2:0] v_9961_0;
  wire [2:0] v_9962_0;
  wire [2:0] v_9963_0;
  wire [2:0] v_9964_0;
  wire [2:0] v_9965_0;
  wire [2:0] v_9966_0;
  wire [2:0] v_9967_0;
  wire [2:0] v_9968_0;
  wire [2:0] v_9969_0;
  wire [2:0] v_9970_0;
  wire [2:0] v_9971_0;
  wire [2:0] v_9972_0;
  wire [2:0] v_9973_0;
  wire [2:0] v_9974_0;
  wire [2:0] v_9975_0;
  wire [2:0] v_9976_0;
  wire [2:0] v_9977_0;
  wire [2:0] v_9978_0;
  wire [2:0] v_9979_0;
  wire [2:0] v_9980_0;
  wire [2:0] v_9981_0;
  wire [2:0] v_9982_0;
  wire [2:0] v_9983_0;
  wire [2:0] v_9984_0;
  wire [2:0] v_9985_0;
  wire [2:0] v_9986_0;
  wire [2:0] v_9987_0;
  wire [2:0] v_9988_0;
  wire [2:0] v_9989_0;
  wire [2:0] v_9990_0;
  wire [2:0] v_9991_0;
  wire [2:0] v_9992_0;
  wire [2:0] v_9993_0;
  wire [2:0] v_9994_0;
  wire [2:0] v_9995_0;
  wire [2:0] v_9996_0;
  wire [2:0] v_9997_0;
  wire [2:0] v_9998_0;
  wire [2:0] v_9999_0;
  wire [2:0] v_10000_0;
  wire [2:0] v_10001_0;
  wire [2:0] v_10002_0;
  wire [2:0] v_10003_0;
  wire [2:0] v_10004_0;
  wire [2:0] v_10005_0;
  wire [2:0] v_10006_0;
  wire [2:0] v_10007_0;
  wire [2:0] v_10008_0;
  wire [2:0] v_10009_0;
  wire [2:0] v_10010_0;
  wire [2:0] v_10011_0;
  wire [2:0] v_10012_0;
  wire [2:0] v_10013_0;
  wire [2:0] v_10014_0;
  wire [2:0] v_10015_0;
  wire [2:0] v_10016_0;
  wire [2:0] v_10017_0;
  wire [2:0] v_10018_0;
  wire [2:0] v_10019_0;
  wire [2:0] v_10020_0;
  wire [2:0] v_10021_0;
  wire [2:0] v_10022_0;
  wire [2:0] v_10023_0;
  wire [2:0] v_10024_0;
  wire [2:0] v_10025_0;
  wire [2:0] v_10026_0;
  wire [2:0] v_10027_0;
  wire [2:0] v_10028_0;
  wire [2:0] v_10029_0;
  wire [2:0] v_10030_0;
  wire [2:0] v_10031_0;
  wire [2:0] v_10032_0;
  wire [2:0] v_10033_0;
  wire [2:0] v_10034_0;
  wire [2:0] v_10035_0;
  wire [2:0] v_10036_0;
  wire [2:0] v_10037_0;
  wire [2:0] v_10038_0;
  wire [2:0] v_10039_0;
  wire [2:0] v_10040_0;
  wire [2:0] v_10041_0;
  wire [2:0] v_10042_0;
  wire [2:0] v_10043_0;
  wire [2:0] v_10044_0;
  wire [2:0] v_10045_0;
  wire [2:0] v_10046_0;
  wire [2:0] v_10047_0;
  wire [2:0] v_10048_0;
  wire [2:0] v_10049_0;
  wire [2:0] v_10050_0;
  wire [2:0] v_10051_0;
  wire [2:0] v_10052_0;
  wire [2:0] v_10053_0;
  wire [2:0] v_10054_0;
  wire [2:0] v_10055_0;
  wire [2:0] v_10056_0;
  wire [2:0] v_10057_0;
  wire [2:0] v_10058_0;
  wire [2:0] v_10059_0;
  wire [2:0] v_10060_0;
  wire [2:0] v_10061_0;
  wire [2:0] v_10062_0;
  wire [2:0] v_10063_0;
  wire [2:0] v_10064_0;
  wire [2:0] v_10065_0;
  wire [2:0] v_10066_0;
  wire [2:0] v_10067_0;
  wire [2:0] v_10068_0;
  wire [2:0] v_10069_0;
  wire [2:0] v_10070_0;
  wire [2:0] v_10071_0;
  wire [2:0] v_10072_0;
  wire [2:0] v_10073_0;
  wire [2:0] v_10074_0;
  wire [2:0] v_10075_0;
  wire [2:0] v_10076_0;
  wire [2:0] v_10077_0;
  wire [2:0] v_10078_0;
  wire [2:0] v_10079_0;
  wire [2:0] v_10080_0;
  wire [2:0] v_10081_0;
  wire [2:0] v_10082_0;
  wire [2:0] v_10083_0;
  wire [2:0] v_10084_0;
  wire [2:0] v_10085_0;
  wire [2:0] v_10086_0;
  wire [2:0] v_10087_0;
  wire [2:0] v_10088_0;
  wire [2:0] v_10089_0;
  wire [2:0] v_10090_0;
  wire [2:0] v_10091_0;
  wire [2:0] v_10092_0;
  wire [2:0] v_10093_0;
  wire [2:0] v_10094_0;
  wire [2:0] v_10095_0;
  wire [2:0] v_10096_0;
  wire [2:0] v_10097_0;
  wire [2:0] v_10098_0;
  wire [2:0] v_10099_0;
  wire [2:0] v_10100_0;
  wire [2:0] v_10101_0;
  wire [2:0] v_10102_0;
  wire [2:0] v_10103_0;
  wire [2:0] v_10104_0;
  wire [2:0] v_10105_0;
  wire [2:0] v_10106_0;
  wire [2:0] v_10107_0;
  wire [2:0] v_10108_0;
  wire [2:0] v_10109_0;
  wire [2:0] v_10110_0;
  wire [2:0] v_10111_0;
  wire [2:0] v_10112_0;
  wire [2:0] v_10113_0;
  wire [2:0] v_10114_0;
  wire [2:0] v_10115_0;
  wire [2:0] v_10116_0;
  wire [2:0] v_10117_0;
  wire [2:0] v_10118_0;
  wire [2:0] v_10119_0;
  wire [2:0] v_10120_0;
  wire [2:0] v_10121_0;
  wire [2:0] v_10122_0;
  wire [2:0] v_10123_0;
  wire [2:0] v_10124_0;
  wire [2:0] v_10125_0;
  wire [2:0] v_10126_0;
  wire [2:0] v_10127_0;
  wire [2:0] v_10128_0;
  wire [2:0] v_10129_0;
  wire [2:0] v_10130_0;
  wire [2:0] v_10131_0;
  wire [2:0] v_10132_0;
  wire [2:0] v_10133_0;
  wire [2:0] v_10134_0;
  wire [2:0] v_10135_0;
  wire [2:0] v_10136_0;
  wire [2:0] v_10137_0;
  wire [2:0] v_10138_0;
  wire [2:0] v_10139_0;
  wire [2:0] v_10140_0;
  wire [2:0] v_10141_0;
  wire [2:0] v_10142_0;
  wire [2:0] v_10143_0;
  wire [2:0] v_10144_0;
  wire [2:0] v_10145_0;
  wire [2:0] v_10146_0;
  wire [2:0] v_10147_0;
  wire [2:0] v_10148_0;
  wire [2:0] v_10149_0;
  wire [2:0] v_10150_0;
  wire [2:0] v_10151_0;
  wire [2:0] v_10152_0;
  wire [2:0] v_10153_0;
  wire [2:0] v_10154_0;
  wire [2:0] v_10155_0;
  wire [2:0] v_10156_0;
  wire [2:0] v_10157_0;
  wire [2:0] v_10158_0;
  wire [2:0] v_10159_0;
  wire [2:0] v_10160_0;
  wire [2:0] v_10161_0;
  wire [2:0] v_10162_0;
  wire [2:0] v_10163_0;
  wire [2:0] v_10164_0;
  wire [2:0] v_10165_0;
  wire [2:0] v_10166_0;
  wire [2:0] v_10167_0;
  wire [2:0] v_10168_0;
  wire [2:0] v_10169_0;
  wire [2:0] v_10170_0;
  wire [2:0] v_10171_0;
  wire [2:0] v_10172_0;
  wire [2:0] v_10173_0;
  wire [2:0] v_10174_0;
  wire [2:0] v_10175_0;
  wire [2:0] v_10176_0;
  wire [2:0] v_10177_0;
  wire [2:0] v_10178_0;
  wire [2:0] v_10179_0;
  wire [2:0] v_10180_0;
  wire [2:0] v_10181_0;
  wire [2:0] v_10182_0;
  wire [2:0] v_10183_0;
  wire [2:0] v_10184_0;
  wire [2:0] v_10185_0;
  wire [2:0] v_10186_0;
  wire [2:0] v_10187_0;
  wire [2:0] v_10188_0;
  wire [2:0] v_10189_0;
  wire [2:0] v_10190_0;
  wire [2:0] v_10191_0;
  wire [2:0] v_10192_0;
  wire [2:0] v_10193_0;
  wire [2:0] v_10194_0;
  wire [2:0] v_10195_0;
  wire [2:0] v_10196_0;
  wire [2:0] v_10197_0;
  wire [2:0] v_10198_0;
  wire [2:0] v_10199_0;
  wire [2:0] v_10200_0;
  wire [2:0] v_10201_0;
  wire [2:0] v_10202_0;
  wire [2:0] v_10203_0;
  wire [2:0] v_10204_0;
  wire [2:0] v_10205_0;
  wire [2:0] v_10206_0;
  wire [2:0] v_10207_0;
  wire [2:0] v_10208_0;
  wire [2:0] v_10209_0;
  wire [2:0] v_10210_0;
  wire [2:0] v_10211_0;
  wire [2:0] v_10212_0;
  wire [2:0] v_10213_0;
  wire [2:0] v_10214_0;
  wire [2:0] v_10215_0;
  wire [2:0] v_10216_0;
  wire [2:0] v_10217_0;
  wire [2:0] v_10218_0;
  wire [2:0] v_10219_0;
  wire [2:0] v_10220_0;
  wire [2:0] v_10221_0;
  wire [2:0] v_10222_0;
  wire [2:0] v_10223_0;
  wire [2:0] v_10224_0;
  wire [2:0] v_10225_0;
  wire [2:0] v_10226_0;
  wire [2:0] v_10227_0;
  wire [2:0] v_10228_0;
  wire [2:0] v_10229_0;
  wire [2:0] v_10230_0;
  wire [2:0] v_10231_0;
  wire [2:0] v_10232_0;
  wire [2:0] v_10233_0;
  wire [2:0] v_10234_0;
  wire [2:0] v_10235_0;
  wire [2:0] v_10236_0;
  wire [2:0] v_10237_0;
  wire [2:0] v_10238_0;
  wire [2:0] v_10239_0;
  wire [2:0] v_10240_0;
  wire [2:0] v_10241_0;
  wire [2:0] v_10242_0;
  wire [2:0] v_10243_0;
  wire [2:0] v_10244_0;
  wire [2:0] v_10245_0;
  wire [2:0] v_10246_0;
  wire [2:0] v_10247_0;
  wire [2:0] v_10248_0;
  wire [2:0] v_10249_0;
  wire [2:0] v_10250_0;
  wire [2:0] v_10251_0;
  wire [2:0] v_10252_0;
  wire [2:0] v_10253_0;
  wire [2:0] v_10254_0;
  wire [2:0] v_10255_0;
  wire [2:0] v_10256_0;
  wire [2:0] v_10257_0;
  wire [2:0] v_10258_0;
  wire [2:0] v_10259_0;
  wire [2:0] v_10260_0;
  wire [2:0] v_10261_0;
  wire [2:0] v_10262_0;
  wire [2:0] v_10263_0;
  wire [2:0] v_10264_0;
  wire [2:0] v_10265_0;
  wire [2:0] v_10266_0;
  wire [2:0] v_10267_0;
  wire [2:0] v_10268_0;
  wire [2:0] v_10269_0;
  wire [2:0] v_10270_0;
  wire [2:0] v_10271_0;
  wire [2:0] v_10272_0;
  wire [2:0] v_10273_0;
  wire [2:0] v_10274_0;
  wire [2:0] v_10275_0;
  wire [2:0] v_10276_0;
  wire [2:0] v_10277_0;
  wire [2:0] v_10278_0;
  wire [2:0] v_10279_0;
  wire [2:0] v_10280_0;
  wire [2:0] v_10281_0;
  wire [2:0] v_10282_0;
  wire [2:0] v_10283_0;
  wire [2:0] v_10284_0;
  wire [2:0] v_10285_0;
  wire [2:0] v_10286_0;
  wire [2:0] v_10287_0;
  wire [2:0] v_10288_0;
  wire [2:0] v_10289_0;
  wire [2:0] v_10290_0;
  wire [2:0] v_10291_0;
  wire [2:0] v_10292_0;
  wire [2:0] v_10293_0;
  wire [2:0] v_10294_0;
  wire [2:0] v_10295_0;
  wire [2:0] v_10296_0;
  wire [2:0] v_10297_0;
  wire [2:0] v_10298_0;
  wire [2:0] v_10299_0;
  wire [2:0] v_10300_0;
  wire [2:0] v_10301_0;
  wire [2:0] v_10302_0;
  wire [2:0] v_10303_0;
  wire [2:0] v_10304_0;
  wire [2:0] v_10305_0;
  wire [2:0] v_10306_0;
  wire [2:0] v_10307_0;
  wire [2:0] v_10308_0;
  wire [2:0] v_10309_0;
  wire [2:0] v_10310_0;
  wire [2:0] v_10311_0;
  wire [2:0] v_10312_0;
  wire [2:0] v_10313_0;
  wire [2:0] v_10314_0;
  wire [2:0] v_10315_0;
  wire [2:0] v_10316_0;
  wire [2:0] v_10317_0;
  wire [2:0] v_10318_0;
  wire [2:0] v_10319_0;
  wire [2:0] v_10320_0;
  wire [2:0] v_10321_0;
  wire [2:0] v_10322_0;
  wire [2:0] v_10323_0;
  wire [2:0] v_10324_0;
  wire [2:0] v_10325_0;
  wire [2:0] v_10326_0;
  wire [2:0] v_10327_0;
  wire [2:0] v_10328_0;
  wire [2:0] v_10329_0;
  wire [2:0] v_10330_0;
  wire [2:0] v_10331_0;
  wire [2:0] v_10332_0;
  wire [2:0] v_10333_0;
  wire [2:0] v_10334_0;
  wire [2:0] v_10335_0;
  wire [2:0] v_10336_0;
  wire [2:0] v_10337_0;
  wire [2:0] v_10338_0;
  wire [2:0] v_10339_0;
  wire [2:0] v_10340_0;
  wire [2:0] v_10341_0;
  wire [2:0] v_10342_0;
  wire [2:0] v_10343_0;
  wire [2:0] v_10344_0;
  wire [2:0] v_10345_0;
  wire [2:0] v_10346_0;
  wire [2:0] v_10347_0;
  wire [2:0] v_10348_0;
  wire [2:0] v_10349_0;
  wire [2:0] v_10350_0;
  wire [2:0] v_10351_0;
  wire [2:0] v_10352_0;
  wire [2:0] v_10353_0;
  wire [2:0] v_10354_0;
  wire [2:0] v_10355_0;
  wire [2:0] v_10356_0;
  wire [2:0] v_10357_0;
  wire [2:0] v_10358_0;
  wire [2:0] v_10359_0;
  wire [2:0] v_10360_0;
  wire [2:0] v_10361_0;
  wire [2:0] v_10362_0;
  wire [2:0] v_10363_0;
  wire [2:0] v_10364_0;
  wire [2:0] v_10365_0;
  wire [2:0] v_10366_0;
  wire [2:0] v_10367_0;
  wire [2:0] v_10368_0;
  wire [2:0] v_10369_0;
  wire [2:0] v_10370_0;
  wire [2:0] v_10371_0;
  wire [2:0] v_10372_0;
  wire [2:0] v_10373_0;
  wire [2:0] v_10374_0;
  wire [2:0] v_10375_0;
  wire [2:0] v_10376_0;
  wire [2:0] v_10377_0;
  wire [2:0] v_10378_0;
  wire [2:0] v_10379_0;
  wire [2:0] v_10380_0;
  wire [2:0] v_10381_0;
  wire [2:0] v_10382_0;
  wire [2:0] v_10383_0;
  wire [2:0] v_10384_0;
  wire [2:0] v_10385_0;
  wire [2:0] v_10386_0;
  wire [2:0] v_10387_0;
  wire [2:0] v_10388_0;
  wire [2:0] v_10389_0;
  wire [2:0] v_10390_0;
  wire [2:0] v_10391_0;
  wire [2:0] v_10392_0;
  wire [2:0] v_10393_0;
  wire [2:0] v_10394_0;
  wire [2:0] v_10395_0;
  wire [2:0] v_10396_0;
  wire [2:0] v_10397_0;
  wire [2:0] v_10398_0;
  wire [2:0] v_10399_0;
  wire [2:0] v_10400_0;
  wire [2:0] v_10401_0;
  wire [2:0] v_10402_0;
  wire [2:0] v_10403_0;
  wire [2:0] v_10404_0;
  wire [2:0] v_10405_0;
  wire [2:0] v_10406_0;
  wire [2:0] v_10407_0;
  wire [2:0] v_10408_0;
  wire [2:0] v_10409_0;
  wire [2:0] v_10410_0;
  wire [2:0] v_10411_0;
  wire [2:0] v_10412_0;
  wire [2:0] v_10413_0;
  wire [2:0] v_10414_0;
  wire [2:0] v_10415_0;
  wire [2:0] v_10416_0;
  wire [2:0] v_10417_0;
  wire [2:0] v_10418_0;
  wire [2:0] v_10419_0;
  wire [2:0] v_10420_0;
  wire [2:0] v_10421_0;
  wire [2:0] v_10422_0;
  wire [2:0] v_10423_0;
  wire [2:0] v_10424_0;
  wire [2:0] v_10425_0;
  wire [2:0] v_10426_0;
  wire [2:0] v_10427_0;
  wire [2:0] v_10428_0;
  wire [2:0] v_10429_0;
  wire [2:0] v_10430_0;
  wire [2:0] v_10431_0;
  wire [2:0] v_10432_0;
  wire [2:0] v_10433_0;
  wire [2:0] v_10434_0;
  wire [2:0] v_10435_0;
  wire [2:0] v_10436_0;
  wire [2:0] v_10437_0;
  wire [2:0] v_10438_0;
  wire [2:0] v_10439_0;
  wire [2:0] v_10440_0;
  wire [2:0] v_10441_0;
  wire [2:0] v_10442_0;
  wire [2:0] v_10443_0;
  wire [2:0] v_10444_0;
  wire [2:0] v_10445_0;
  wire [2:0] v_10446_0;
  wire [2:0] v_10447_0;
  wire [2:0] v_10448_0;
  wire [2:0] v_10449_0;
  wire [2:0] v_10450_0;
  wire [2:0] v_10451_0;
  wire [2:0] v_10452_0;
  wire [2:0] v_10453_0;
  wire [2:0] v_10454_0;
  wire [2:0] v_10455_0;
  wire [2:0] v_10456_0;
  wire [2:0] v_10457_0;
  wire [2:0] v_10458_0;
  wire [2:0] v_10459_0;
  wire [2:0] v_10460_0;
  wire [2:0] v_10461_0;
  wire [2:0] v_10462_0;
  wire [2:0] v_10463_0;
  wire [2:0] v_10464_0;
  wire [2:0] v_10465_0;
  wire [2:0] v_10466_0;
  wire [2:0] v_10467_0;
  wire [2:0] v_10468_0;
  wire [2:0] v_10469_0;
  wire [2:0] v_10470_0;
  wire [2:0] v_10471_0;
  wire [2:0] v_10472_0;
  wire [2:0] v_10473_0;
  wire [2:0] v_10474_0;
  wire [2:0] v_10475_0;
  wire [2:0] v_10476_0;
  wire [2:0] v_10477_0;
  wire [2:0] v_10478_0;
  wire [2:0] v_10479_0;
  wire [2:0] v_10480_0;
  wire [2:0] v_10481_0;
  wire [2:0] v_10482_0;
  wire [2:0] v_10483_0;
  wire [2:0] v_10484_0;
  wire [2:0] v_10485_0;
  wire [2:0] v_10486_0;
  wire [2:0] v_10487_0;
  wire [2:0] v_10488_0;
  wire [2:0] v_10489_0;
  wire [2:0] v_10490_0;
  wire [2:0] v_10491_0;
  wire [2:0] v_10492_0;
  wire [2:0] v_10493_0;
  wire [2:0] v_10494_0;
  wire [2:0] v_10495_0;
  wire [2:0] v_10496_0;
  wire [2:0] v_10497_0;
  wire [2:0] v_10498_0;
  wire [2:0] v_10499_0;
  wire [2:0] v_10500_0;
  wire [2:0] v_10501_0;
  wire [2:0] v_10502_0;
  wire [2:0] v_10503_0;
  wire [2:0] v_10504_0;
  wire [2:0] v_10505_0;
  wire [2:0] v_10506_0;
  wire [2:0] v_10507_0;
  wire [2:0] v_10508_0;
  wire [2:0] v_10509_0;
  wire [2:0] v_10510_0;
  wire [2:0] v_10511_0;
  wire [2:0] v_10512_0;
  wire [2:0] v_10513_0;
  wire [2:0] v_10514_0;
  wire [2:0] v_10515_0;
  wire [2:0] v_10516_0;
  wire [2:0] v_10517_0;
  wire [2:0] v_10518_0;
  wire [2:0] v_10519_0;
  wire [2:0] v_10520_0;
  wire [2:0] v_10521_0;
  wire [2:0] v_10522_0;
  wire [2:0] v_10523_0;
  wire [2:0] v_10524_0;
  wire [2:0] v_10525_0;
  wire [2:0] v_10526_0;
  wire [2:0] v_10527_0;
  wire [2:0] v_10528_0;
  wire [2:0] v_10529_0;
  wire [2:0] v_10530_0;
  wire [2:0] v_10531_0;
  wire [2:0] v_10532_0;
  wire [2:0] v_10533_0;
  wire [2:0] v_10534_0;
  wire [2:0] v_10535_0;
  wire [2:0] v_10536_0;
  wire [2:0] v_10537_0;
  wire [2:0] v_10538_0;
  wire [2:0] v_10539_0;
  wire [2:0] v_10540_0;
  wire [2:0] v_10541_0;
  wire [2:0] v_10542_0;
  wire [2:0] v_10543_0;
  wire [2:0] v_10544_0;
  wire [2:0] v_10545_0;
  wire [2:0] v_10546_0;
  wire [2:0] v_10547_0;
  wire [2:0] v_10548_0;
  wire [2:0] v_10549_0;
  wire [2:0] v_10550_0;
  wire [2:0] v_10551_0;
  wire [2:0] v_10552_0;
  wire [2:0] v_10553_0;
  wire [2:0] v_10554_0;
  wire [2:0] v_10555_0;
  wire [2:0] v_10556_0;
  wire [2:0] v_10557_0;
  wire [2:0] v_10558_0;
  wire [2:0] v_10559_0;
  wire [2:0] v_10560_0;
  wire [2:0] v_10561_0;
  wire [2:0] v_10562_0;
  wire [2:0] v_10563_0;
  wire [2:0] v_10564_0;
  wire [2:0] v_10565_0;
  wire [2:0] v_10566_0;
  wire [2:0] v_10567_0;
  wire [2:0] v_10568_0;
  wire [2:0] v_10569_0;
  wire [2:0] v_10570_0;
  wire [2:0] v_10571_0;
  wire [2:0] v_10572_0;
  wire [2:0] v_10573_0;
  wire [2:0] v_10574_0;
  wire [2:0] v_10575_0;
  wire [2:0] v_10576_0;
  wire [2:0] v_10577_0;
  wire [2:0] v_10578_0;
  wire [2:0] v_10579_0;
  wire [2:0] v_10580_0;
  wire [2:0] v_10581_0;
  wire [2:0] v_10582_0;
  wire [2:0] v_10583_0;
  wire [2:0] v_10584_0;
  wire [2:0] v_10585_0;
  wire [2:0] v_10586_0;
  wire [2:0] v_10587_0;
  wire [2:0] v_10588_0;
  wire [2:0] v_10589_0;
  wire [2:0] v_10590_0;
  wire [2:0] v_10591_0;
  wire [2:0] v_10592_0;
  wire [2:0] v_10593_0;
  wire [2:0] v_10594_0;
  wire [2:0] v_10595_0;
  wire [2:0] v_10596_0;
  wire [2:0] v_10597_0;
  wire [2:0] v_10598_0;
  wire [2:0] v_10599_0;
  wire [2:0] v_10600_0;
  wire [2:0] v_10601_0;
  wire [2:0] v_10602_0;
  wire [2:0] v_10603_0;
  wire [2:0] v_10604_0;
  wire [2:0] v_10605_0;
  wire [2:0] v_10606_0;
  wire [2:0] v_10607_0;
  wire [2:0] v_10608_0;
  wire [2:0] v_10609_0;
  wire [2:0] v_10610_0;
  wire [2:0] v_10611_0;
  wire [2:0] v_10612_0;
  wire [2:0] v_10613_0;
  wire [2:0] v_10614_0;
  wire [2:0] v_10615_0;
  wire [2:0] v_10616_0;
  wire [2:0] v_10617_0;
  wire [2:0] v_10618_0;
  wire [2:0] v_10619_0;
  wire [2:0] v_10620_0;
  wire [2:0] v_10621_0;
  wire [2:0] v_10622_0;
  wire [2:0] v_10623_0;
  wire [2:0] v_10624_0;
  wire [2:0] v_10625_0;
  wire [2:0] v_10626_0;
  wire [2:0] v_10627_0;
  wire [2:0] v_10628_0;
  wire [2:0] v_10629_0;
  wire [2:0] v_10630_0;
  wire [2:0] v_10631_0;
  wire [2:0] v_10632_0;
  wire [2:0] v_10633_0;
  wire [2:0] v_10634_0;
  wire [2:0] v_10635_0;
  wire [2:0] v_10636_0;
  wire [2:0] v_10637_0;
  wire [2:0] v_10638_0;
  wire [2:0] v_10639_0;
  wire [2:0] v_10640_0;
  wire [2:0] v_10641_0;
  wire [2:0] v_10642_0;
  wire [2:0] v_10643_0;
  wire [2:0] v_10644_0;
  wire [2:0] v_10645_0;
  wire [2:0] v_10646_0;
  wire [2:0] v_10647_0;
  wire [2:0] v_10648_0;
  wire [2:0] v_10649_0;
  wire [2:0] v_10650_0;
  wire [2:0] v_10651_0;
  wire [2:0] v_10652_0;
  wire [2:0] v_10653_0;
  wire [2:0] v_10654_0;
  wire [2:0] v_10655_0;
  wire [2:0] v_10656_0;
  wire [2:0] v_10657_0;
  wire [2:0] v_10658_0;
  wire [2:0] v_10659_0;
  wire [2:0] v_10660_0;
  wire [2:0] v_10661_0;
  wire [2:0] v_10662_0;
  wire [2:0] v_10663_0;
  wire [2:0] v_10664_0;
  wire [2:0] v_10665_0;
  wire [2:0] v_10666_0;
  wire [2:0] v_10667_0;
  wire [2:0] v_10668_0;
  wire [2:0] v_10669_0;
  wire [2:0] v_10670_0;
  wire [2:0] v_10671_0;
  wire [2:0] v_10672_0;
  wire [2:0] v_10673_0;
  wire [2:0] v_10674_0;
  wire [2:0] v_10675_0;
  wire [2:0] v_10676_0;
  wire [2:0] v_10677_0;
  wire [2:0] v_10678_0;
  wire [2:0] v_10679_0;
  wire [2:0] v_10680_0;
  wire [2:0] v_10681_0;
  wire [2:0] v_10682_0;
  wire [2:0] v_10683_0;
  wire [2:0] v_10684_0;
  wire [2:0] v_10685_0;
  wire [2:0] v_10686_0;
  wire [2:0] v_10687_0;
  wire [2:0] v_10688_0;
  wire [2:0] v_10689_0;
  wire [2:0] v_10690_0;
  wire [2:0] v_10691_0;
  wire [2:0] v_10692_0;
  wire [2:0] v_10693_0;
  wire [2:0] v_10694_0;
  wire [2:0] v_10695_0;
  wire [2:0] v_10696_0;
  wire [2:0] v_10697_0;
  wire [2:0] v_10698_0;
  wire [2:0] v_10699_0;
  wire [2:0] v_10700_0;
  wire [2:0] v_10701_0;
  wire [2:0] v_10702_0;
  wire [2:0] v_10703_0;
  wire [2:0] v_10704_0;
  wire [2:0] v_10705_0;
  wire [2:0] v_10706_0;
  wire [2:0] v_10707_0;
  wire [2:0] v_10708_0;
  wire [2:0] v_10709_0;
  wire [2:0] v_10710_0;
  wire [2:0] v_10711_0;
  wire [2:0] v_10712_0;
  wire [2:0] v_10713_0;
  wire [2:0] v_10714_0;
  wire [2:0] v_10715_0;
  wire [2:0] v_10716_0;
  wire [2:0] v_10717_0;
  wire [2:0] v_10718_0;
  wire [2:0] v_10719_0;
  wire [2:0] v_10720_0;
  wire [2:0] v_10721_0;
  wire [2:0] v_10722_0;
  wire [2:0] v_10723_0;
  wire [2:0] v_10724_0;
  wire [2:0] v_10725_0;
  wire [2:0] v_10726_0;
  wire [2:0] v_10727_0;
  wire [2:0] v_10728_0;
  wire [2:0] v_10729_0;
  wire [2:0] v_10730_0;
  wire [2:0] v_10731_0;
  wire [2:0] v_10732_0;
  wire [2:0] v_10733_0;
  wire [2:0] v_10734_0;
  wire [2:0] v_10735_0;
  wire [2:0] v_10736_0;
  wire [2:0] v_10737_0;
  wire [2:0] v_10738_0;
  wire [2:0] v_10739_0;
  wire [2:0] v_10740_0;
  wire [2:0] v_10741_0;
  wire [2:0] v_10742_0;
  wire [2:0] v_10743_0;
  wire [2:0] v_10744_0;
  wire [2:0] v_10745_0;
  wire [2:0] v_10746_0;
  wire [2:0] v_10747_0;
  wire [2:0] v_10748_0;
  wire [2:0] v_10749_0;
  wire [2:0] v_10750_0;
  wire [2:0] v_10751_0;
  wire [2:0] v_10752_0;
  wire [2:0] v_10753_0;
  wire [2:0] v_10754_0;
  wire [2:0] v_10755_0;
  wire [2:0] v_10756_0;
  wire [2:0] v_10757_0;
  wire [2:0] v_10758_0;
  wire [2:0] v_10759_0;
  wire [2:0] v_10760_0;
  wire [2:0] v_10761_0;
  wire [2:0] v_10762_0;
  wire [2:0] v_10763_0;
  wire [2:0] v_10764_0;
  wire [2:0] v_10765_0;
  wire [2:0] v_10766_0;
  wire [2:0] v_10767_0;
  wire [2:0] v_10768_0;
  wire [2:0] v_10769_0;
  wire [2:0] v_10770_0;
  wire [2:0] v_10771_0;
  wire [2:0] v_10772_0;
  wire [2:0] v_10773_0;
  wire [2:0] v_10774_0;
  wire [2:0] v_10775_0;
  wire [2:0] v_10776_0;
  wire [2:0] v_10777_0;
  wire [2:0] v_10778_0;
  wire [2:0] v_10779_0;
  wire [2:0] v_10780_0;
  wire [2:0] v_10781_0;
  wire [2:0] v_10782_0;
  wire [2:0] v_10783_0;
  wire [2:0] v_10784_0;
  wire [2:0] v_10785_0;
  wire [2:0] v_10786_0;
  wire [2:0] v_10787_0;
  wire [2:0] v_10788_0;
  wire [2:0] v_10789_0;
  wire [2:0] v_10790_0;
  wire [2:0] v_10791_0;
  wire [2:0] v_10792_0;
  wire [2:0] v_10793_0;
  wire [2:0] v_10794_0;
  wire [2:0] v_10795_0;
  wire [2:0] v_10796_0;
  wire [2:0] v_10797_0;
  wire [2:0] v_10798_0;
  wire [2:0] v_10799_0;
  wire [2:0] v_10800_0;
  wire [2:0] v_10801_0;
  wire [2:0] v_10802_0;
  wire [2:0] v_10803_0;
  wire [2:0] v_10804_0;
  wire [2:0] v_10805_0;
  wire [2:0] v_10806_0;
  wire [2:0] v_10807_0;
  wire [2:0] v_10808_0;
  wire [2:0] v_10809_0;
  wire [2:0] v_10810_0;
  wire [2:0] v_10811_0;
  wire [2:0] v_10812_0;
  wire [2:0] v_10813_0;
  wire [2:0] v_10814_0;
  wire [2:0] v_10815_0;
  wire [2:0] v_10816_0;
  wire [2:0] v_10817_0;
  wire [2:0] v_10818_0;
  wire [2:0] v_10819_0;
  wire [2:0] v_10820_0;
  wire [2:0] v_10821_0;
  wire [2:0] v_10822_0;
  wire [2:0] v_10823_0;
  wire [2:0] v_10824_0;
  wire [2:0] v_10825_0;
  wire [2:0] v_10826_0;
  wire [2:0] v_10827_0;
  wire [2:0] v_10828_0;
  wire [2:0] v_10829_0;
  wire [2:0] v_10830_0;
  wire [2:0] v_10831_0;
  wire [2:0] v_10832_0;
  wire [2:0] v_10833_0;
  wire [2:0] v_10834_0;
  wire [2:0] v_10835_0;
  wire [2:0] v_10836_0;
  wire [2:0] v_10837_0;
  wire [2:0] v_10838_0;
  wire [2:0] v_10839_0;
  wire [2:0] v_10840_0;
  wire [2:0] v_10841_0;
  wire [2:0] v_10842_0;
  wire [2:0] v_10843_0;
  wire [2:0] v_10844_0;
  wire [2:0] v_10845_0;
  wire [2:0] v_10846_0;
  wire [2:0] v_10847_0;
  wire [2:0] v_10848_0;
  wire [2:0] v_10849_0;
  wire [2:0] v_10850_0;
  wire [2:0] v_10851_0;
  wire [2:0] v_10852_0;
  wire [2:0] v_10853_0;
  wire [2:0] v_10854_0;
  wire [2:0] v_10855_0;
  wire [2:0] v_10856_0;
  wire [2:0] v_10857_0;
  wire [2:0] v_10858_0;
  wire [2:0] v_10859_0;
  wire [2:0] v_10860_0;
  wire [2:0] v_10861_0;
  wire [2:0] v_10862_0;
  wire [2:0] v_10863_0;
  wire [2:0] v_10864_0;
  wire [2:0] v_10865_0;
  wire [2:0] v_10866_0;
  wire [2:0] v_10867_0;
  wire [2:0] v_10868_0;
  wire [2:0] v_10869_0;
  wire [2:0] v_10870_0;
  wire [2:0] v_10871_0;
  wire [2:0] v_10872_0;
  wire [2:0] v_10873_0;
  wire [2:0] v_10874_0;
  wire [2:0] v_10875_0;
  wire [2:0] v_10876_0;
  wire [2:0] v_10877_0;
  wire [2:0] v_10878_0;
  wire [2:0] v_10879_0;
  wire [2:0] v_10880_0;
  wire [2:0] v_10881_0;
  wire [2:0] v_10882_0;
  wire [2:0] v_10883_0;
  wire [2:0] v_10884_0;
  wire [2:0] v_10885_0;
  wire [2:0] v_10886_0;
  wire [2:0] v_10887_0;
  wire [2:0] v_10888_0;
  wire [2:0] v_10889_0;
  wire [2:0] v_10890_0;
  wire [2:0] v_10891_0;
  wire [2:0] v_10892_0;
  wire [2:0] v_10893_0;
  wire [2:0] v_10894_0;
  wire [2:0] v_10895_0;
  wire [2:0] v_10896_0;
  wire [2:0] v_10897_0;
  wire [2:0] v_10898_0;
  wire [2:0] v_10899_0;
  wire [2:0] v_10900_0;
  wire [2:0] v_10901_0;
  wire [2:0] v_10902_0;
  wire [2:0] v_10903_0;
  wire [2:0] v_10904_0;
  wire [2:0] v_10905_0;
  wire [2:0] v_10906_0;
  wire [2:0] v_10907_0;
  wire [2:0] v_10908_0;
  wire [2:0] v_10909_0;
  wire [2:0] v_10910_0;
  wire [2:0] v_10911_0;
  wire [2:0] v_10912_0;
  wire [2:0] v_10913_0;
  wire [2:0] v_10914_0;
  wire [2:0] v_10915_0;
  wire [2:0] v_10916_0;
  wire [2:0] v_10917_0;
  wire [2:0] v_10918_0;
  wire [2:0] v_10919_0;
  wire [2:0] v_10920_0;
  wire [2:0] v_10921_0;
  wire [2:0] v_10922_0;
  wire [2:0] v_10923_0;
  wire [2:0] v_10924_0;
  wire [2:0] v_10925_0;
  wire [2:0] v_10926_0;
  wire [2:0] v_10927_0;
  wire [2:0] v_10928_0;
  wire [2:0] v_10929_0;
  wire [2:0] v_10930_0;
  wire [2:0] v_10931_0;
  wire [2:0] v_10932_0;
  wire [2:0] v_10933_0;
  wire [2:0] v_10934_0;
  wire [2:0] v_10935_0;
  wire [2:0] v_10936_0;
  wire [2:0] v_10937_0;
  wire [2:0] v_10938_0;
  wire [2:0] v_10939_0;
  wire [2:0] v_10940_0;
  wire [2:0] v_10941_0;
  wire [2:0] v_10942_0;
  wire [2:0] v_10943_0;
  wire [2:0] v_10944_0;
  wire [2:0] v_10945_0;
  wire [2:0] v_10946_0;
  wire [2:0] v_10947_0;
  wire [2:0] v_10948_0;
  wire [2:0] v_10949_0;
  wire [2:0] v_10950_0;
  wire [2:0] v_10951_0;
  wire [2:0] v_10952_0;
  wire [2:0] v_10953_0;
  wire [2:0] v_10954_0;
  wire [2:0] v_10955_0;
  wire [2:0] v_10956_0;
  wire [2:0] v_10957_0;
  wire [2:0] v_10958_0;
  wire [2:0] v_10959_0;
  wire [2:0] v_10960_0;
  wire [2:0] v_10961_0;
  wire [2:0] v_10962_0;
  wire [2:0] v_10963_0;
  wire [2:0] v_10964_0;
  wire [2:0] v_10965_0;
  wire [2:0] v_10966_0;
  wire [2:0] v_10967_0;
  wire [2:0] v_10968_0;
  wire [2:0] v_10969_0;
  wire [2:0] v_10970_0;
  wire [2:0] v_10971_0;
  wire [2:0] v_10972_0;
  wire [2:0] v_10973_0;
  wire [2:0] v_10974_0;
  wire [2:0] v_10975_0;
  wire [2:0] v_10976_0;
  wire [2:0] v_10977_0;
  wire [2:0] v_10978_0;
  wire [2:0] v_10979_0;
  wire [2:0] v_10980_0;
  wire [2:0] v_10981_0;
  wire [2:0] v_10982_0;
  wire [2:0] v_10983_0;
  wire [2:0] v_10984_0;
  wire [2:0] v_10985_0;
  wire [2:0] v_10986_0;
  wire [2:0] v_10987_0;
  wire [2:0] v_10988_0;
  wire [2:0] v_10989_0;
  wire [2:0] v_10990_0;
  wire [2:0] v_10991_0;
  wire [2:0] v_10992_0;
  wire [2:0] v_10993_0;
  wire [2:0] v_10994_0;
  wire [2:0] v_10995_0;
  wire [2:0] v_10996_0;
  wire [2:0] v_10997_0;
  wire [2:0] v_10998_0;
  wire [2:0] v_10999_0;
  wire [2:0] v_11000_0;
  wire [2:0] v_11001_0;
  wire [2:0] v_11002_0;
  wire [2:0] v_11003_0;
  wire [2:0] v_11004_0;
  wire [2:0] v_11005_0;
  wire [2:0] v_11006_0;
  wire [2:0] v_11007_0;
  wire [2:0] v_11008_0;
  wire [2:0] v_11009_0;
  wire [2:0] v_11010_0;
  wire [2:0] v_11011_0;
  wire [2:0] v_11012_0;
  wire [2:0] v_11013_0;
  wire [2:0] v_11014_0;
  wire [2:0] v_11015_0;
  wire [2:0] v_11016_0;
  wire [2:0] v_11017_0;
  wire [2:0] v_11018_0;
  wire [2:0] v_11019_0;
  wire [2:0] v_11020_0;
  wire [2:0] v_11021_0;
  wire [2:0] v_11022_0;
  wire [2:0] v_11023_0;
  wire [2:0] v_11024_0;
  wire [2:0] v_11025_0;
  wire [2:0] v_11026_0;
  wire [2:0] v_11027_0;
  wire [2:0] v_11028_0;
  wire [2:0] v_11029_0;
  wire [2:0] v_11030_0;
  wire [2:0] v_11031_0;
  wire [2:0] v_11032_0;
  wire [2:0] v_11033_0;
  wire [2:0] v_11034_0;
  wire [2:0] v_11035_0;
  wire [2:0] v_11036_0;
  wire [2:0] v_11037_0;
  wire [2:0] v_11038_0;
  wire [2:0] v_11039_0;
  wire [2:0] v_11040_0;
  wire [2:0] v_11041_0;
  wire [2:0] v_11042_0;
  wire [2:0] v_11043_0;
  wire [2:0] v_11044_0;
  wire [2:0] v_11045_0;
  wire [2:0] v_11046_0;
  wire [2:0] v_11047_0;
  wire [2:0] v_11048_0;
  wire [2:0] v_11049_0;
  wire [2:0] v_11050_0;
  wire [2:0] v_11051_0;
  wire [2:0] v_11052_0;
  wire [2:0] v_11053_0;
  wire [2:0] v_11054_0;
  wire [2:0] v_11055_0;
  wire [2:0] v_11056_0;
  wire [2:0] v_11057_0;
  wire [2:0] v_11058_0;
  wire [2:0] v_11059_0;
  wire [2:0] v_11060_0;
  wire [2:0] v_11061_0;
  wire [2:0] v_11062_0;
  wire [2:0] v_11063_0;
  wire [2:0] v_11064_0;
  wire [2:0] v_11065_0;
  wire [2:0] v_11066_0;
  wire [2:0] v_11067_0;
  wire [2:0] v_11068_0;
  wire [2:0] v_11069_0;
  wire [2:0] v_11070_0;
  wire [2:0] v_11071_0;
  wire [2:0] v_11072_0;
  wire [2:0] v_11073_0;
  wire [2:0] v_11074_0;
  wire [2:0] v_11075_0;
  wire [2:0] v_11076_0;
  wire [2:0] v_11077_0;
  wire [2:0] v_11078_0;
  wire [2:0] v_11079_0;
  wire [2:0] v_11080_0;
  wire [2:0] v_11081_0;
  wire [2:0] v_11082_0;
  wire [2:0] v_11083_0;
  wire [2:0] v_11084_0;
  wire [2:0] v_11085_0;
  wire [2:0] v_11086_0;
  wire [2:0] v_11087_0;
  wire [2:0] v_11088_0;
  wire [2:0] v_11089_0;
  wire [2:0] v_11090_0;
  wire [2:0] v_11091_0;
  wire [2:0] v_11092_0;
  wire [2:0] v_11093_0;
  wire [2:0] v_11094_0;
  wire [2:0] v_11095_0;
  wire [2:0] v_11096_0;
  wire [2:0] v_11097_0;
  wire [2:0] v_11098_0;
  wire [2:0] v_11099_0;
  wire [2:0] v_11100_0;
  wire [2:0] v_11101_0;
  wire [2:0] v_11102_0;
  wire [2:0] v_11103_0;
  wire [2:0] v_11104_0;
  wire [2:0] v_11105_0;
  wire [2:0] v_11106_0;
  wire [2:0] v_11107_0;
  wire [2:0] v_11108_0;
  wire [2:0] v_11109_0;
  wire [2:0] v_11110_0;
  wire [2:0] v_11111_0;
  wire [2:0] v_11112_0;
  wire [2:0] v_11113_0;
  wire [2:0] v_11114_0;
  wire [2:0] v_11115_0;
  wire [2:0] v_11116_0;
  wire [2:0] v_11117_0;
  wire [2:0] v_11118_0;
  wire [2:0] v_11119_0;
  wire [2:0] v_11120_0;
  wire [2:0] v_11121_0;
  wire [2:0] v_11122_0;
  wire [2:0] v_11123_0;
  wire [2:0] v_11124_0;
  wire [2:0] v_11125_0;
  wire [2:0] v_11126_0;
  wire [2:0] v_11127_0;
  wire [2:0] v_11128_0;
  wire [2:0] v_11129_0;
  wire [2:0] v_11130_0;
  wire [2:0] v_11131_0;
  wire [2:0] v_11132_0;
  wire [2:0] v_11133_0;
  wire [2:0] v_11134_0;
  wire [2:0] v_11135_0;
  wire [2:0] v_11136_0;
  wire [2:0] v_11137_0;
  wire [2:0] v_11138_0;
  wire [2:0] v_11139_0;
  wire [2:0] v_11140_0;
  wire [2:0] v_11141_0;
  wire [2:0] v_11142_0;
  wire [2:0] v_11143_0;
  wire [2:0] v_11144_0;
  wire [2:0] v_11145_0;
  wire [2:0] v_11146_0;
  wire [2:0] v_11147_0;
  wire [2:0] v_11148_0;
  wire [2:0] v_11149_0;
  wire [2:0] v_11150_0;
  wire [2:0] v_11151_0;
  wire [2:0] v_11152_0;
  wire [2:0] v_11153_0;
  wire [2:0] v_11154_0;
  wire [2:0] v_11155_0;
  wire [2:0] v_11156_0;
  wire [2:0] v_11157_0;
  wire [2:0] v_11158_0;
  wire [2:0] v_11159_0;
  wire [2:0] v_11160_0;
  wire [2:0] v_11161_0;
  wire [2:0] v_11162_0;
  wire [2:0] v_11163_0;
  wire [2:0] v_11164_0;
  wire [2:0] v_11165_0;
  wire [2:0] v_11166_0;
  wire [2:0] v_11167_0;
  wire [2:0] v_11168_0;
  wire [2:0] v_11169_0;
  wire [2:0] v_11170_0;
  wire [2:0] v_11171_0;
  wire [2:0] v_11172_0;
  wire [2:0] v_11173_0;
  wire [2:0] v_11174_0;
  wire [2:0] v_11175_0;
  wire [2:0] v_11176_0;
  wire [2:0] v_11177_0;
  wire [2:0] v_11178_0;
  wire [2:0] v_11179_0;
  wire [2:0] v_11180_0;
  wire [2:0] v_11181_0;
  wire [2:0] v_11182_0;
  wire [2:0] v_11183_0;
  wire [2:0] v_11184_0;
  wire [2:0] v_11185_0;
  wire [2:0] v_11186_0;
  wire [2:0] v_11187_0;
  wire [2:0] v_11188_0;
  wire [2:0] v_11189_0;
  wire [2:0] v_11190_0;
  wire [2:0] v_11191_0;
  wire [2:0] v_11192_0;
  wire [2:0] v_11193_0;
  wire [2:0] v_11194_0;
  wire [2:0] v_11195_0;
  wire [2:0] v_11196_0;
  wire [2:0] v_11197_0;
  wire [2:0] v_11198_0;
  wire [2:0] v_11199_0;
  wire [2:0] v_11200_0;
  wire [2:0] v_11201_0;
  wire [2:0] v_11202_0;
  wire [2:0] v_11203_0;
  wire [2:0] v_11204_0;
  wire [2:0] v_11205_0;
  wire [2:0] v_11206_0;
  wire [2:0] v_11207_0;
  wire [2:0] v_11208_0;
  wire [2:0] v_11209_0;
  wire [2:0] v_11210_0;
  wire [2:0] v_11211_0;
  wire [2:0] v_11212_0;
  wire [2:0] v_11213_0;
  wire [2:0] v_11214_0;
  wire [2:0] v_11215_0;
  wire [2:0] v_11216_0;
  wire [2:0] v_11217_0;
  wire [2:0] v_11218_0;
  wire [2:0] v_11219_0;
  wire [2:0] v_11220_0;
  wire [2:0] v_11221_0;
  wire [2:0] v_11222_0;
  wire [2:0] v_11223_0;
  wire [2:0] v_11224_0;
  wire [2:0] v_11225_0;
  wire [2:0] v_11226_0;
  wire [2:0] v_11227_0;
  wire [2:0] v_11228_0;
  wire [2:0] v_11229_0;
  wire [2:0] v_11230_0;
  wire [2:0] v_11231_0;
  wire [2:0] v_11232_0;
  wire [2:0] v_11233_0;
  wire [2:0] v_11234_0;
  wire [2:0] v_11235_0;
  wire [2:0] v_11236_0;
  wire [2:0] v_11237_0;
  wire [2:0] v_11238_0;
  wire [2:0] v_11239_0;
  wire [2:0] v_11240_0;
  wire [2:0] v_11241_0;
  wire [2:0] v_11242_0;
  wire [2:0] v_11243_0;
  wire [2:0] v_11244_0;
  wire [2:0] v_11245_0;
  wire [2:0] v_11246_0;
  wire [2:0] v_11247_0;
  wire [2:0] v_11248_0;
  wire [2:0] v_11249_0;
  wire [2:0] v_11250_0;
  wire [2:0] v_11251_0;
  wire [2:0] v_11252_0;
  wire [2:0] v_11253_0;
  wire [2:0] v_11254_0;
  wire [2:0] v_11255_0;
  wire [2:0] v_11256_0;
  wire [2:0] v_11257_0;
  wire [2:0] v_11258_0;
  wire [2:0] v_11259_0;
  wire [2:0] v_11260_0;
  wire [2:0] v_11261_0;
  wire [2:0] v_11262_0;
  wire [2:0] v_11263_0;
  wire [2:0] v_11264_0;
  wire [2:0] v_11265_0;
  wire [2:0] v_11266_0;
  wire [2:0] v_11267_0;
  wire [2:0] v_11268_0;
  wire [2:0] v_11269_0;
  wire [2:0] v_11270_0;
  wire [2:0] v_11271_0;
  wire [2:0] v_11272_0;
  wire [2:0] v_11273_0;
  wire [2:0] v_11274_0;
  wire [2:0] v_11275_0;
  wire [2:0] v_11276_0;
  wire [2:0] v_11277_0;
  wire [2:0] v_11278_0;
  wire [2:0] v_11279_0;
  wire [2:0] v_11280_0;
  wire [2:0] v_11281_0;
  wire [2:0] v_11282_0;
  wire [2:0] v_11283_0;
  wire [2:0] v_11284_0;
  wire [2:0] v_11285_0;
  wire [2:0] v_11286_0;
  wire [2:0] v_11287_0;
  wire [2:0] v_11288_0;
  wire [2:0] v_11289_0;
  wire [2:0] v_11290_0;
  wire [2:0] v_11291_0;
  wire [2:0] v_11292_0;
  wire [2:0] v_11293_0;
  wire [2:0] v_11294_0;
  wire [2:0] v_11295_0;
  wire [2:0] v_11296_0;
  wire [2:0] v_11297_0;
  wire [2:0] v_11298_0;
  wire [2:0] v_11299_0;
  wire [2:0] v_11300_0;
  wire [2:0] v_11301_0;
  wire [2:0] v_11302_0;
  wire [2:0] v_11303_0;
  wire [2:0] v_11304_0;
  wire [2:0] v_11305_0;
  wire [2:0] v_11306_0;
  wire [2:0] v_11307_0;
  wire [2:0] v_11308_0;
  wire [2:0] v_11309_0;
  wire [2:0] v_11310_0;
  wire [2:0] v_11311_0;
  wire [2:0] v_11312_0;
  wire [2:0] v_11313_0;
  wire [2:0] v_11314_0;
  wire [2:0] v_11315_0;
  wire [2:0] v_11316_0;
  wire [2:0] v_11317_0;
  wire [2:0] v_11318_0;
  wire [2:0] v_11319_0;
  wire [2:0] v_11320_0;
  wire [2:0] v_11321_0;
  wire [2:0] v_11322_0;
  wire [2:0] v_11323_0;
  wire [2:0] v_11324_0;
  wire [2:0] v_11325_0;
  wire [2:0] v_11326_0;
  wire [2:0] v_11327_0;
  wire [2:0] v_11328_0;
  wire [2:0] v_11329_0;
  wire [2:0] v_11330_0;
  wire [2:0] v_11331_0;
  wire [2:0] v_11332_0;
  wire [2:0] v_11333_0;
  wire [2:0] v_11334_0;
  wire [2:0] v_11335_0;
  wire [2:0] v_11336_0;
  wire [2:0] v_11337_0;
  wire [2:0] v_11338_0;
  wire [2:0] v_11339_0;
  wire [2:0] v_11340_0;
  wire [2:0] v_11341_0;
  wire [2:0] v_11342_0;
  wire [2:0] v_11343_0;
  wire [2:0] v_11344_0;
  wire [2:0] v_11345_0;
  wire [2:0] v_11346_0;
  wire [2:0] v_11347_0;
  wire [2:0] v_11348_0;
  wire [2:0] v_11349_0;
  wire [2:0] v_11350_0;
  wire [2:0] v_11351_0;
  wire [2:0] v_11352_0;
  wire [2:0] v_11353_0;
  wire [2:0] v_11354_0;
  wire [2:0] v_11355_0;
  wire [2:0] v_11356_0;
  wire [2:0] v_11357_0;
  wire [2:0] v_11358_0;
  wire [2:0] v_11359_0;
  wire [2:0] v_11360_0;
  wire [2:0] v_11361_0;
  wire [2:0] v_11362_0;
  wire [2:0] v_11363_0;
  wire [2:0] v_11364_0;
  wire [2:0] v_11365_0;
  wire [2:0] v_11366_0;
  wire [2:0] v_11367_0;
  wire [2:0] v_11368_0;
  wire [2:0] v_11369_0;
  wire [2:0] v_11370_0;
  wire [2:0] v_11371_0;
  wire [2:0] v_11372_0;
  wire [2:0] v_11373_0;
  wire [2:0] v_11374_0;
  wire [2:0] v_11375_0;
  wire [2:0] v_11376_0;
  wire [2:0] v_11377_0;
  wire [2:0] v_11378_0;
  wire [2:0] v_11379_0;
  wire [2:0] v_11380_0;
  wire [2:0] v_11381_0;
  wire [2:0] v_11382_0;
  wire [2:0] v_11383_0;
  wire [2:0] v_11384_0;
  wire [2:0] v_11385_0;
  wire [2:0] v_11386_0;
  wire [2:0] v_11387_0;
  wire [2:0] v_11388_0;
  wire [2:0] v_11389_0;
  wire [2:0] v_11390_0;
  wire [2:0] v_11391_0;
  wire [2:0] v_11392_0;
  wire [2:0] v_11393_0;
  wire [2:0] v_11394_0;
  wire [2:0] v_11395_0;
  wire [2:0] v_11396_0;
  wire [2:0] v_11397_0;
  wire [2:0] v_11398_0;
  wire [2:0] v_11399_0;
  wire [2:0] v_11400_0;
  wire [2:0] v_11401_0;
  wire [2:0] v_11402_0;
  wire [2:0] v_11403_0;
  wire [2:0] v_11404_0;
  wire [2:0] v_11405_0;
  wire [2:0] v_11406_0;
  wire [2:0] v_11407_0;
  wire [2:0] v_11408_0;
  wire [2:0] v_11409_0;
  wire [2:0] v_11410_0;
  wire [2:0] v_11411_0;
  wire [2:0] v_11412_0;
  wire [2:0] v_11413_0;
  wire [2:0] v_11414_0;
  wire [2:0] v_11415_0;
  wire [2:0] v_11416_0;
  wire [2:0] v_11417_0;
  wire [2:0] v_11418_0;
  wire [2:0] v_11419_0;
  wire [2:0] v_11420_0;
  wire [2:0] v_11421_0;
  wire [2:0] v_11422_0;
  wire [2:0] v_11423_0;
  wire [2:0] v_11424_0;
  wire [2:0] v_11425_0;
  wire [2:0] v_11426_0;
  wire [2:0] v_11427_0;
  wire [2:0] v_11428_0;
  wire [2:0] v_11429_0;
  wire [2:0] v_11430_0;
  wire [2:0] v_11431_0;
  wire [2:0] v_11432_0;
  wire [2:0] v_11433_0;
  wire [2:0] v_11434_0;
  wire [2:0] v_11435_0;
  wire [2:0] v_11436_0;
  wire [2:0] v_11437_0;
  wire [2:0] v_11438_0;
  wire [2:0] v_11439_0;
  wire [2:0] v_11440_0;
  wire [2:0] v_11441_0;
  wire [2:0] v_11442_0;
  wire [2:0] v_11443_0;
  wire [2:0] v_11444_0;
  wire [2:0] v_11445_0;
  wire [2:0] v_11446_0;
  wire [2:0] v_11447_0;
  wire [2:0] v_11448_0;
  wire [2:0] v_11449_0;
  wire [2:0] v_11450_0;
  wire [2:0] v_11451_0;
  wire [2:0] v_11452_0;
  wire [2:0] v_11453_0;
  wire [2:0] v_11454_0;
  wire [2:0] v_11455_0;
  wire [2:0] v_11456_0;
  wire [2:0] v_11457_0;
  wire [2:0] v_11458_0;
  wire [2:0] v_11459_0;
  wire [2:0] v_11460_0;
  wire [2:0] v_11461_0;
  wire [2:0] v_11462_0;
  wire [2:0] v_11463_0;
  wire [2:0] v_11464_0;
  wire [2:0] v_11465_0;
  wire [2:0] v_11466_0;
  wire [2:0] v_11467_0;
  wire [2:0] v_11468_0;
  wire [2:0] v_11469_0;
  wire [2:0] v_11470_0;
  wire [2:0] v_11471_0;
  wire [2:0] v_11472_0;
  wire [2:0] v_11473_0;
  wire [2:0] v_11474_0;
  wire [2:0] v_11475_0;
  wire [2:0] v_11476_0;
  wire [2:0] v_11477_0;
  wire [2:0] v_11478_0;
  wire [2:0] v_11479_0;
  wire [2:0] v_11480_0;
  wire [2:0] v_11481_0;
  wire [2:0] v_11482_0;
  wire [2:0] v_11483_0;
  wire [2:0] v_11484_0;
  wire [2:0] v_11485_0;
  wire [2:0] v_11486_0;
  wire [2:0] v_11487_0;
  wire [2:0] v_11488_0;
  wire [2:0] v_11489_0;
  wire [2:0] v_11490_0;
  wire [2:0] v_11491_0;
  wire [2:0] v_11492_0;
  wire [2:0] v_11493_0;
  wire [2:0] v_11494_0;
  wire [2:0] v_11495_0;
  wire [2:0] v_11496_0;
  wire [2:0] v_11497_0;
  wire [2:0] v_11498_0;
  wire [2:0] v_11499_0;
  wire [2:0] v_11500_0;
  wire [2:0] v_11501_0;
  wire [2:0] v_11502_0;
  wire [2:0] v_11503_0;
  wire [2:0] v_11504_0;
  wire [2:0] v_11505_0;
  wire [2:0] v_11506_0;
  wire [2:0] v_11507_0;
  wire [2:0] v_11508_0;
  wire [2:0] v_11509_0;
  wire [2:0] v_11510_0;
  wire [2:0] v_11511_0;
  wire [2:0] v_11512_0;
  wire [2:0] v_11513_0;
  wire [2:0] v_11514_0;
  wire [2:0] v_11515_0;
  wire [2:0] v_11516_0;
  wire [2:0] v_11517_0;
  wire [2:0] v_11518_0;
  wire [2:0] v_11519_0;
  wire [2:0] v_11520_0;
  wire [2:0] v_11521_0;
  wire [2:0] v_11522_0;
  wire [2:0] v_11523_0;
  wire [2:0] v_11524_0;
  wire [2:0] v_11525_0;
  wire [2:0] v_11526_0;
  wire [2:0] v_11527_0;
  wire [2:0] v_11528_0;
  wire [2:0] v_11529_0;
  wire [2:0] v_11530_0;
  wire [2:0] v_11531_0;
  wire [2:0] v_11532_0;
  wire [2:0] v_11533_0;
  wire [2:0] v_11534_0;
  wire [2:0] v_11535_0;
  wire [2:0] v_11536_0;
  wire [2:0] v_11537_0;
  wire [2:0] v_11538_0;
  wire [2:0] v_11539_0;
  wire [2:0] v_11540_0;
  wire [2:0] v_11541_0;
  wire [2:0] v_11542_0;
  wire [2:0] v_11543_0;
  wire [2:0] v_11544_0;
  wire [2:0] v_11545_0;
  wire [2:0] v_11546_0;
  wire [2:0] v_11547_0;
  wire [2:0] v_11548_0;
  wire [2:0] v_11549_0;
  wire [2:0] v_11550_0;
  wire [2:0] v_11551_0;
  wire [2:0] v_11552_0;
  wire [2:0] v_11553_0;
  wire [2:0] v_11554_0;
  wire [2:0] v_11555_0;
  wire [2:0] v_11556_0;
  wire [2:0] v_11557_0;
  wire [2:0] v_11558_0;
  wire [2:0] v_11559_0;
  wire [2:0] v_11560_0;
  wire [2:0] v_11561_0;
  wire [2:0] v_11562_0;
  wire [2:0] v_11563_0;
  wire [2:0] v_11564_0;
  wire [2:0] v_11565_0;
  wire [2:0] v_11566_0;
  wire [2:0] v_11567_0;
  wire [2:0] v_11568_0;
  wire [2:0] v_11569_0;
  wire [2:0] v_11570_0;
  wire [2:0] v_11571_0;
  wire [2:0] v_11572_0;
  wire [2:0] v_11573_0;
  wire [2:0] v_11574_0;
  wire [2:0] v_11575_0;
  wire [2:0] v_11576_0;
  wire [2:0] v_11577_0;
  wire [2:0] v_11578_0;
  wire [2:0] v_11579_0;
  wire [2:0] v_11580_0;
  wire [2:0] v_11581_0;
  wire [2:0] v_11582_0;
  wire [2:0] v_11583_0;
  wire [2:0] v_11584_0;
  wire [2:0] v_11585_0;
  wire [2:0] v_11586_0;
  wire [2:0] v_11587_0;
  wire [2:0] v_11588_0;
  wire [2:0] v_11589_0;
  wire [2:0] v_11590_0;
  wire [2:0] v_11591_0;
  wire [2:0] v_11592_0;
  wire [2:0] v_11593_0;
  wire [2:0] v_11594_0;
  wire [2:0] v_11595_0;
  wire [2:0] v_11596_0;
  wire [2:0] v_11597_0;
  wire [2:0] v_11598_0;
  wire [2:0] v_11599_0;
  wire [2:0] v_11600_0;
  wire [2:0] v_11601_0;
  wire [2:0] v_11602_0;
  wire [2:0] v_11603_0;
  wire [2:0] v_11604_0;
  wire [2:0] v_11605_0;
  wire [2:0] v_11606_0;
  wire [2:0] v_11607_0;
  wire [2:0] v_11608_0;
  wire [2:0] v_11609_0;
  wire [2:0] v_11610_0;
  wire [2:0] v_11611_0;
  wire [2:0] v_11612_0;
  wire [2:0] v_11613_0;
  wire [2:0] v_11614_0;
  wire [2:0] v_11615_0;
  wire [2:0] v_11616_0;
  wire [2:0] v_11617_0;
  wire [2:0] v_11618_0;
  wire [2:0] v_11619_0;
  wire [2:0] v_11620_0;
  wire [2:0] v_11621_0;
  wire [2:0] v_11622_0;
  wire [2:0] v_11623_0;
  wire [2:0] v_11624_0;
  wire [2:0] v_11625_0;
  wire [2:0] v_11626_0;
  wire [2:0] v_11627_0;
  wire [2:0] v_11628_0;
  wire [2:0] v_11629_0;
  wire [2:0] v_11630_0;
  wire [2:0] v_11631_0;
  wire [2:0] v_11632_0;
  wire [2:0] v_11633_0;
  wire [2:0] v_11634_0;
  wire [2:0] v_11635_0;
  wire [2:0] v_11636_0;
  wire [2:0] v_11637_0;
  wire [2:0] v_11638_0;
  wire [2:0] v_11639_0;
  wire [2:0] v_11640_0;
  wire [2:0] v_11641_0;
  wire [2:0] v_11642_0;
  wire [2:0] v_11643_0;
  wire [2:0] v_11644_0;
  wire [2:0] v_11645_0;
  wire [2:0] v_11646_0;
  wire [2:0] v_11647_0;
  wire [2:0] v_11648_0;
  wire [2:0] v_11649_0;
  wire [2:0] v_11650_0;
  wire [2:0] v_11651_0;
  wire [2:0] v_11652_0;
  wire [2:0] v_11653_0;
  wire [2:0] v_11654_0;
  wire [2:0] v_11655_0;
  wire [2:0] v_11656_0;
  wire [2:0] v_11657_0;
  wire [2:0] v_11658_0;
  wire [2:0] v_11659_0;
  wire [2:0] v_11660_0;
  wire [2:0] v_11661_0;
  wire [2:0] v_11662_0;
  wire [2:0] v_11663_0;
  wire [2:0] v_11664_0;
  wire [2:0] v_11665_0;
  wire [2:0] v_11666_0;
  wire [2:0] v_11667_0;
  wire [2:0] v_11668_0;
  wire [2:0] v_11669_0;
  wire [2:0] v_11670_0;
  wire [2:0] v_11671_0;
  wire [2:0] v_11672_0;
  wire [2:0] v_11673_0;
  wire [2:0] v_11674_0;
  wire [2:0] v_11675_0;
  wire [2:0] v_11676_0;
  wire [2:0] v_11677_0;
  wire [2:0] v_11678_0;
  wire [2:0] v_11679_0;
  wire [2:0] v_11680_0;
  wire [2:0] v_11681_0;
  wire [2:0] v_11682_0;
  wire [2:0] v_11683_0;
  wire [2:0] v_11684_0;
  wire [2:0] v_11685_0;
  wire [2:0] v_11686_0;
  wire [2:0] v_11687_0;
  wire [2:0] v_11688_0;
  wire [2:0] v_11689_0;
  wire [2:0] v_11690_0;
  wire [2:0] v_11691_0;
  wire [2:0] v_11692_0;
  wire [2:0] v_11693_0;
  wire [2:0] v_11694_0;
  wire [2:0] v_11695_0;
  wire [2:0] v_11696_0;
  wire [2:0] v_11697_0;
  wire [2:0] v_11698_0;
  wire [2:0] v_11699_0;
  wire [2:0] v_11700_0;
  wire [2:0] v_11701_0;
  wire [2:0] v_11702_0;
  wire [2:0] v_11703_0;
  wire [2:0] v_11704_0;
  wire [2:0] v_11705_0;
  wire [2:0] v_11706_0;
  wire [2:0] v_11707_0;
  wire [2:0] v_11708_0;
  wire [2:0] v_11709_0;
  wire [2:0] v_11710_0;
  wire [2:0] v_11711_0;
  wire [2:0] v_11712_0;
  wire [2:0] v_11713_0;
  wire [2:0] v_11714_0;
  wire [2:0] v_11715_0;
  wire [2:0] v_11716_0;
  wire [2:0] v_11717_0;
  wire [2:0] v_11718_0;
  wire [2:0] v_11719_0;
  wire [2:0] v_11720_0;
  wire [2:0] v_11721_0;
  wire [2:0] v_11722_0;
  wire [2:0] v_11723_0;
  wire [2:0] v_11724_0;
  wire [2:0] v_11725_0;
  wire [2:0] v_11726_0;
  wire [2:0] v_11727_0;
  wire [2:0] v_11728_0;
  wire [2:0] v_11729_0;
  wire [2:0] v_11730_0;
  wire [2:0] v_11731_0;
  wire [2:0] v_11732_0;
  wire [2:0] v_11733_0;
  wire [2:0] v_11734_0;
  wire [2:0] v_11735_0;
  wire [2:0] v_11736_0;
  wire [2:0] v_11737_0;
  wire [2:0] v_11738_0;
  wire [2:0] v_11739_0;
  wire [2:0] v_11740_0;
  wire [2:0] v_11741_0;
  wire [2:0] v_11742_0;
  wire [2:0] v_11743_0;
  wire [2:0] v_11744_0;
  wire [2:0] v_11745_0;
  wire [2:0] v_11746_0;
  wire [2:0] v_11747_0;
  wire [2:0] v_11748_0;
  wire [2:0] v_11749_0;
  wire [2:0] v_11750_0;
  wire [2:0] v_11751_0;
  wire [2:0] v_11752_0;
  wire [2:0] v_11753_0;
  wire [2:0] v_11754_0;
  wire [2:0] v_11755_0;
  wire [2:0] v_11756_0;
  wire [2:0] v_11757_0;
  wire [2:0] v_11758_0;
  wire [2:0] v_11759_0;
  wire [2:0] v_11760_0;
  wire [2:0] v_11761_0;
  wire [2:0] v_11762_0;
  wire [2:0] v_11763_0;
  wire [2:0] v_11764_0;
  wire [2:0] v_11765_0;
  wire [2:0] v_11766_0;
  wire [2:0] v_11767_0;
  wire [2:0] v_11768_0;
  wire [2:0] v_11769_0;
  wire [2:0] v_11770_0;
  wire [2:0] v_11771_0;
  wire [2:0] v_11772_0;
  wire [2:0] v_11773_0;
  wire [2:0] v_11774_0;
  wire [2:0] v_11775_0;
  wire [2:0] v_11776_0;
  wire [2:0] v_11777_0;
  wire [2:0] v_11778_0;
  wire [2:0] v_11779_0;
  wire [2:0] v_11780_0;
  wire [2:0] v_11781_0;
  wire [2:0] v_11782_0;
  wire [2:0] v_11783_0;
  wire [2:0] v_11784_0;
  wire [2:0] v_11785_0;
  wire [2:0] v_11786_0;
  wire [2:0] v_11787_0;
  wire [2:0] v_11788_0;
  wire [2:0] v_11789_0;
  wire [2:0] v_11790_0;
  wire [2:0] v_11791_0;
  wire [2:0] v_11792_0;
  wire [2:0] v_11793_0;
  wire [2:0] v_11794_0;
  wire [2:0] v_11795_0;
  wire [2:0] v_11796_0;
  wire [2:0] v_11797_0;
  wire [2:0] v_11798_0;
  wire [2:0] v_11799_0;
  wire [2:0] v_11800_0;
  wire [2:0] v_11801_0;
  wire [2:0] v_11802_0;
  wire [2:0] v_11803_0;
  wire [2:0] v_11804_0;
  wire [2:0] v_11805_0;
  wire [2:0] v_11806_0;
  wire [2:0] v_11807_0;
  wire [2:0] v_11808_0;
  wire [2:0] v_11809_0;
  wire [2:0] v_11810_0;
  wire [2:0] v_11811_0;
  wire [2:0] v_11812_0;
  wire [2:0] v_11813_0;
  wire [2:0] v_11814_0;
  wire [2:0] v_11815_0;
  wire [2:0] v_11816_0;
  wire [2:0] v_11817_0;
  wire [2:0] v_11818_0;
  wire [2:0] v_11819_0;
  wire [2:0] v_11820_0;
  wire [2:0] v_11821_0;
  wire [2:0] v_11822_0;
  wire [2:0] v_11823_0;
  wire [2:0] v_11824_0;
  wire [2:0] v_11825_0;
  wire [2:0] v_11826_0;
  wire [2:0] v_11827_0;
  wire [2:0] v_11828_0;
  wire [2:0] v_11829_0;
  wire [2:0] v_11830_0;
  wire [2:0] v_11831_0;
  wire [2:0] v_11832_0;
  wire [2:0] v_11833_0;
  wire [2:0] v_11834_0;
  wire [2:0] v_11835_0;
  wire [2:0] v_11836_0;
  wire [2:0] v_11837_0;
  wire [2:0] v_11838_0;
  wire [2:0] v_11839_0;
  wire [2:0] v_11840_0;
  wire [2:0] v_11841_0;
  wire [2:0] v_11842_0;
  wire [2:0] v_11843_0;
  wire [2:0] v_11844_0;
  wire [2:0] v_11845_0;
  wire [2:0] v_11846_0;
  wire [2:0] v_11847_0;
  wire [2:0] v_11848_0;
  wire [2:0] v_11849_0;
  wire [2:0] v_11850_0;
  wire [2:0] v_11851_0;
  wire [2:0] v_11852_0;
  wire [2:0] v_11853_0;
  wire [2:0] v_11854_0;
  wire [2:0] v_11855_0;
  wire [2:0] v_11856_0;
  wire [2:0] v_11857_0;
  wire [2:0] v_11858_0;
  wire [2:0] v_11859_0;
  wire [2:0] v_11860_0;
  wire [2:0] v_11861_0;
  wire [2:0] v_11862_0;
  wire [2:0] v_11863_0;
  wire [2:0] v_11864_0;
  wire [2:0] v_11865_0;
  wire [2:0] v_11866_0;
  wire [2:0] v_11867_0;
  wire [2:0] v_11868_0;
  wire [2:0] v_11869_0;
  wire [2:0] v_11870_0;
  wire [2:0] v_11871_0;
  wire [2:0] v_11872_0;
  wire [2:0] v_11873_0;
  wire [2:0] v_11874_0;
  wire [2:0] v_11875_0;
  wire [2:0] v_11876_0;
  wire [2:0] v_11877_0;
  wire [2:0] v_11878_0;
  wire [2:0] v_11879_0;
  wire [2:0] v_11880_0;
  wire [2:0] v_11881_0;
  wire [2:0] v_11882_0;
  wire [2:0] v_11883_0;
  wire [2:0] v_11884_0;
  wire [2:0] v_11885_0;
  wire [2:0] v_11886_0;
  wire [2:0] v_11887_0;
  wire [2:0] v_11888_0;
  wire [2:0] v_11889_0;
  wire [2:0] v_11890_0;
  wire [2:0] v_11891_0;
  wire [2:0] v_11892_0;
  wire [2:0] v_11893_0;
  wire [2:0] v_11894_0;
  wire [2:0] v_11895_0;
  wire [2:0] v_11896_0;
  wire [2:0] v_11897_0;
  wire [2:0] v_11898_0;
  wire [2:0] v_11899_0;
  wire [2:0] v_11900_0;
  wire [2:0] v_11901_0;
  wire [2:0] v_11902_0;
  wire [2:0] v_11903_0;
  wire [2:0] v_11904_0;
  wire [2:0] v_11905_0;
  wire [2:0] v_11906_0;
  wire [2:0] v_11907_0;
  wire [2:0] v_11908_0;
  wire [2:0] v_11909_0;
  wire [2:0] v_11910_0;
  wire [2:0] v_11911_0;
  wire [2:0] v_11912_0;
  wire [2:0] v_11913_0;
  wire [2:0] v_11914_0;
  wire [2:0] v_11915_0;
  wire [2:0] v_11916_0;
  wire [2:0] v_11917_0;
  wire [2:0] v_11918_0;
  wire [2:0] v_11919_0;
  wire [2:0] v_11920_0;
  wire [2:0] v_11921_0;
  wire [2:0] v_11922_0;
  wire [2:0] v_11923_0;
  wire [2:0] v_11924_0;
  wire [2:0] v_11925_0;
  wire [2:0] v_11926_0;
  wire [2:0] v_11927_0;
  wire [2:0] v_11928_0;
  wire [2:0] v_11929_0;
  wire [2:0] v_11930_0;
  wire [2:0] v_11931_0;
  wire [2:0] v_11932_0;
  wire [2:0] v_11933_0;
  wire [2:0] v_11934_0;
  wire [2:0] v_11935_0;
  wire [2:0] v_11936_0;
  wire [2:0] v_11937_0;
  wire [2:0] v_11938_0;
  wire [2:0] v_11939_0;
  wire [2:0] v_11940_0;
  wire [2:0] v_11941_0;
  wire [2:0] v_11942_0;
  wire [2:0] v_11943_0;
  wire [2:0] v_11944_0;
  wire [2:0] v_11945_0;
  wire [2:0] v_11946_0;
  wire [2:0] v_11947_0;
  reg [2:0] v_11948_0 = 3'h0;
  wire [0:0] v_11949_0;
  wire [0:0] v_11950_0;
  wire [0:0] v_11951_0;
  wire [0:0] v_11952_0;
  wire [0:0] v_11953_0;
  wire [2:0] v_11954_0;
  wire [2:0] v_11955_0;
  wire [2:0] v_11956_0;
  wire [2:0] v_11957_0;
  wire [0:0] v_11958_0;
  wire [0:0] v_11959_0;
  reg [0:0] v_11960_0 = 1'h0;
  reg [0:0] v_11961_0 = 1'h0;
  wire [0:0] _act_11962_0;
  wire [0:0] v_11963_0;
  wire [0:0] v_11964_0;
  reg [9:0] v_11965_0 = 10'h0;
  wire [9:0] v_11966_0;
  wire [9:0] v_11967_0;
  wire [9:0] v_11968_0;
  wire [0:0] _act_11969_0;
  wire [0:0] v_11970_0;
  wire [0:0] v_11971_0;
  wire [0:0] v_11972_0;
  wire [0:0] v_11973_0;
  wire [9:0] v_11974_0;
  wire [9:0] v_11975_0;
  wire [9:0] v_11976_0;
  wire [0:0] v_11977_0;
  wire [9:0] v_11978_0;
  wire [9:0] v_11979_0;
  wire [9:0] v_11980_0;
  wire [9:0] v_11981_0;
  wire [9:0] v_11982_0;
  wire [9:0] v_11983_0;
  wire [9:0] v_11984_0;
  wire [9:0] v_11985_0;
  wire [9:0] v_11986_0;
  wire [9:0] v_11987_0;
  wire [9:0] v_11988_0;
  reg [9:0] v_11989_0 = 10'h0;
  wire [0:0] v_11990_0;
  wire [9:0] v_11991_0;
  wire [0:0] v_11992_0;
  reg [9:0] v_11993_0 = 10'h0;
  wire [9:0] v_11994_0;
  wire [9:0] v_11995_0;
  wire [9:0] v_11996_0;
  wire [9:0] v_11997_0;
  wire [9:0] v_11998_0;
  wire [9:0] v_11999_0;
  wire [9:0] v_12000_0;
  wire [0:0] v_12001_0;
  reg [2:0] v_12002_0 = 3'h0;
  wire [2:0] v_12003_0;
  wire [2:0] v_12004_0;
  wire [2:0] v_12005_0;
  wire [2:0] v_12006_0;
  wire [2:0] v_12007_0;
  wire [2:0] v_12008_0;
  wire [2:0] v_12009_0;
  wire [0:0] v_12010_0;
  wire [0:0] v_12011_0;
  wire [0:0] v_12012_0;
  wire [2:0] v_12013_0;
  wire [2:0] v_12013_1;
  wire [9:0] v_12014_0;
  wire [9:0] v_12015_0;
  wire [9:0] v_12016_0;
  wire [0:0] v_12017_0;
  wire [2:0] v_12018_0;
  wire [0:0] v_12019_0;
  wire [0:0] v_12020_0;
  wire [0:0] v_12021_0;
  wire [9:0] v_12022_0;
  wire [9:0] v_12023_0;
  wire [9:0] v_12024_0;
  wire [9:0] v_12025_0;
  wire [9:0] v_12026_0;
  wire [9:0] v_12027_0;
  wire [9:0] v_12028_0;
  wire [0:0] v_12029_0;
  wire [0:0] v_12030_0;
  wire [0:0] v_12031_0;
  wire [2:0] v_12032_0;
  wire [2:0] v_12033_0;
  wire [2:0] v_12034_0;
  wire [2:0] v_12035_0;
  wire [2:0] v_12036_0;
  wire [2:0] v_12037_0;
  wire [2:0] v_12038_0;
  wire [0:0] v_12039_0;
  wire [0:0] v_12040_0;
  wire [0:0] v_12041_0;
  wire [0:0] v_12042_0;
  wire [0:0] v_12043_0;
  wire [0:0] v_12044_0;
  wire [0:0] v_12045_0;
  wire [0:0] v_12046_0;
  wire [0:0] v_12047_0;
  wire [0:0] v_12048_0;
  wire [0:0] v_12049_0;
  wire [0:0] v_12050_0;
  wire [0:0] v_12051_0;
  wire [2:0] v_12052_0;
  wire [2:0] v_12053_0;
  wire [2:0] v_12054_0;
  wire [2:0] v_12055_0;
  wire [2:0] v_12056_0;
  wire [2:0] v_12057_0;
  wire [2:0] v_12058_0;
  wire [2:0] v_12059_0;
  wire [0:0] v_12060_0;
  wire [0:0] v_12061_0;
  wire [0:0] v_12062_0;
  wire [0:0] v_12063_0;
  wire [0:0] v_12064_0;
  reg [0:0] v_12065_0 = 1'h1;
  wire [0:0] v_12066_0;
  wire [0:0] v_12067_0;
  wire [0:0] v_12068_0;
  wire [0:0] v_12069_0;
  wire [0:0] v_12070_0;
  wire [0:0] v_12071_0;
  wire [0:0] v_12072_0;
  wire [0:0] v_12073_0;
  wire [0:0] v_12074_0;
  wire [0:0] v_12075_0;
  wire [0:0] v_12076_0;
  wire [0:0] v_12077_0;
  reg [0:0] v_12078_0 = 1'h0;
  wire [0:0] v_12079_0;
  wire [0:0] v_12080_0;
  wire [0:0] v_12081_0;
  wire [0:0] v_12082_0;
  wire [0:0] v_12083_0;
  wire [0:0] v_12084_0;
  wire [15:0] v_12085_0;
  reg [15:0] v_12086_0 = 16'h0;
  wire [0:0] v_12087_0;
  wire [0:0] v_12088_0;
  wire [0:0] v_12089_0;
  reg [0:0] v_12090_0 = 1'h0;
  wire [0:0] v_12091_0;
  reg [0:0] v_12092_0 = 1'h0;
  wire [0:0] v_12093_0;
  wire [0:0] v_12094_0;
  wire [0:0] _act_12095_0;
  wire [0:0] v_12096_0;
  wire [0:0] v_12097_0;
  wire [0:0] v_12098_0;
  reg [0:0] v_12099_0 = 1'h1;
  wire [0:0] v_12100_0;
  wire [0:0] v_12101_0;
  wire [0:0] v_12102_0;
  wire [4:0] v_12103_0;
  wire [0:0] v_12104_0;
  wire [0:0] v_12105_0;
  wire [0:0] v_12106_0;
  wire [0:0] v_12107_0;
  wire [4:0] v_12108_0;
  reg [4:0] v_12109_0 = 5'h0;
  reg [4:0] v_12110_0 = 5'h0;
  wire [0:0] _act_12111_0;
  wire [0:0] _act_12112_0;
  wire [0:0] v_12113_0;
  wire [0:0] v_12114_0;
  wire [0:0] v_12115_0;
  wire [0:0] v_12116_0;
  wire [0:0] v_12117_0;
  wire [0:0] v_12118_0;
  wire [0:0] v_12119_0;
  wire [0:0] v_12120_0;
  wire [0:0] v_12121_0;
  wire [0:0] v_12122_0;
  wire [0:0] v_12123_0;
  wire [0:0] v_12124_0;
  wire [0:0] v_12125_0;
  wire [0:0] v_12126_0;
  wire [0:0] v_12127_0;
  wire [0:0] v_12128_0;
  wire [0:0] v_12129_0;
  wire [0:0] v_12130_0;
  wire [4:0] v_12131_0;
  wire [0:0] v_12132_0;
  wire [0:0] v_12133_0;
  wire [0:0] v_12134_0;
  wire [0:0] v_12135_0;
  wire [0:0] v_12136_0;
  wire [0:0] v_12137_0;
  wire [0:0] v_12138_0;
  wire [0:0] v_12139_0;
  wire [0:0] v_12140_0;
  wire [0:0] v_12141_0;
  wire [0:0] v_12142_0;
  wire [0:0] v_12143_0;
  wire [0:0] v_12144_0;
  wire [0:0] v_12145_0;
  wire [0:0] v_12146_0;
  wire [0:0] v_12147_0;
  wire [0:0] v_12148_0;
  wire [0:0] v_12149_0;
  wire [0:0] v_12150_0;
  wire [0:0] v_12151_0;
  wire [0:0] v_12152_0;
  wire [0:0] v_12153_0;
  wire [0:0] v_12154_0;
  wire [15:0] v_12155_0;
  reg [15:0] v_12156_0 = 16'h0;
  wire [0:0] v_12157_0;
  wire [0:0] v_12158_0;
  wire [0:0] v_12159_0;
  wire [0:0] v_12160_0;
  wire [0:0] v_12161_0;
  wire [0:0] v_12162_0;
  wire [0:0] v_12163_0;
  wire [0:0] v_12164_0;
  wire [15:0] v_12165_0;
  wire [15:0] v_12166_0;
  wire [15:0] v_12167_0;
  wire [0:0] v_12168_0;
  wire [0:0] v_12169_0;
  reg [0:0] v_12170_0 = 1'h0;
  reg [0:0] v_12171_0 = 1'h0;
  wire [0:0] v_12172_0;
  reg [4:0] v_12173_0 = 5'h0;
  wire [4:0] v_12174_0;
  wire [4:0] v_12175_0;
  wire [4:0] v_12176_0;
  wire [0:0] v_12177_0;
  reg [4:0] v_12178_0 = 5'h0;
  wire [4:0] v_12179_0;
  wire [4:0] v_12180_0;
  wire [4:0] v_12181_0;
  wire [0:0] v_12182_0;
  reg [15:0] v_12183_0 = 16'h0;
  wire [15:0] v_12184_0;
  wire [15:0] v_12185_0;
  wire [15:0] v_12186_0;
  wire [15:0] v_12187_0;
  wire [15:0] v_12188_0;
  wire [0:0] v_12189_0;
  wire [15:0] v_12190_0;
  wire [15:0] v_12191_0;
  wire [15:0] v_12192_0;
  wire [15:0] v_12193_0;
  wire [15:0] v_12194_0;
  wire [15:0] v_12195_0;
  wire [15:0] v_12196_0;
  wire [15:0] v_12197_0;
  wire [15:0] v_12198_0;
  wire [15:0] v_12199_0;
  wire [15:0] v_12200_0;
  wire [15:0] v_12201_0;
  wire [0:0] v_12202_0;
  wire [15:0] v_12203_0;
  wire [15:0] v_12203_1;
  wire [4:0] v_12204_0;
  wire [4:0] v_12205_0;
  wire [4:0] v_12206_0;
  wire [0:0] v_12207_0;
  wire [15:0] v_12208_0;
  wire [0:0] v_12209_0;
  wire [0:0] v_12210_0;
  wire [0:0] v_12211_0;
  wire [4:0] v_12212_0;
  wire [4:0] v_12213_0;
  wire [4:0] v_12214_0;
  wire [0:0] v_12215_0;
  wire [15:0] v_12216_0;
  wire [15:0] v_12217_0;
  wire [15:0] v_12218_0;
  wire [0:0] v_12219_0;
  wire [0:0] v_12220_0;
  wire [0:0] v_12221_0;
  wire [0:0] v_12222_0;
  wire [0:0] v_12223_0;
  wire [15:0] v_12224_0;
  wire [0:0] v_12225_0;
  reg [15:0] v_12226_0 = 16'h0;
  wire [0:0] v_12227_0;
  wire [0:0] v_12228_0;
  wire [0:0] v_12229_0;
  wire [0:0] v_12230_0;
  wire [0:0] v_12231_0;
  wire [0:0] v_12232_0;
  wire [0:0] v_12233_0;
  wire [0:0] v_12234_0;
  wire [0:0] v_12235_0;
  wire [0:0] v_12236_0;
  wire [0:0] v_12237_0;
  wire [0:0] v_12238_0;
  wire [0:0] v_12239_0;
  wire [0:0] v_12240_0;
  wire [0:0] v_12241_0;
  wire [0:0] v_12242_0;
  wire [0:0] v_12243_0;
  wire [15:0] v_12244_0;
  wire [15:0] v_12245_0;
  wire [15:0] v_12246_0;
  wire [15:0] v_12247_0;
  wire [15:0] v_12248_0;
  wire [15:0] v_12249_0;
  wire [15:0] v_12250_0;
  wire [15:0] v_12251_0;
  wire [15:0] v_12252_0;
  wire [15:0] v_12253_0;
  wire [15:0] v_12254_0;
  wire [0:0] v_12255_0;
  wire [0:0] v_12256_0;
  wire [0:0] v_12257_0;
  wire [0:0] v_12258_0;
  wire [0:0] v_12259_0;
  wire [0:0] v_12260_0;
  wire [0:0] v_12261_0;
  wire [0:0] v_12262_0;
  wire [0:0] v_12263_0;
  wire [0:0] v_12264_0;
  wire [0:0] v_12265_0;
  wire [0:0] v_12266_0;
  wire [0:0] v_12268_0;
  wire [0:0] v_12270_0;
  wire [0:0] v_12272_0;
  wire [0:0] v_12273_0;
  wire [0:0] v_12274_0;
  wire [0:0] v_12276_0;
  wire [0:0] v_12278_0;
  wire [0:0] v_12279_0;
  wire [0:0] v_12280_0;
  wire [0:0] v_12282_0;
  wire [0:0] v_12284_0;
  wire [0:0] v_12286_0;
  wire [0:0] v_12287_0;
  reg [0:0] v_12288_0 = 1'h0;
  wire [15:0] v_12289_0;
  wire [0:0] v_12290_0;
  wire [0:0] v_12292_0;
  reg [31:0] v_12294_0 = 32'h0;
  wire [31:0] v_12295_0;
  wire [0:0] v_12297_0;
  wire [0:0] v_12299_0;
  wire [0:0] v_12300_0;
  wire [0:0] v_12301_0;
  wire [0:0] v_12303_0;
  wire [0:0] v_12305_0;
  wire [0:0] v_12307_0;
  wire [0:0] v_12308_0;
  wire [0:0] v_12309_0;
  wire [0:0] v_12311_0;
  wire [0:0] v_12313_0;
  wire [0:0] v_12314_0;
  wire [0:0] v_12315_0;
  wire [0:0] v_12317_0;
  wire [0:0] v_12319_0;
  wire [0:0] v_12322_0;
  wire [0:0] v_12324_0;
  wire [0:0] v_12325_0;
  wire [0:0] v_12327_0;
  wire [0:0] v_12328_0;
  wire [0:0] v_12329_0;
  wire [0:0] v_12330_0;
  wire [0:0] v_12331_0;
  wire [0:0] v_12332_0;
  reg [0:0] v_12334_0 = 1'h0;
  wire [0:0] v_12335_0;
  wire [0:0] v_12336_0;
  wire [0:0] v_12337_0;
  wire [0:0] v_12338_0;
  wire [0:0] v_12339_0;
  wire [0:0] v_12340_0;
  wire [0:0] v_12341_0;
  wire [0:0] v_12342_0;
  wire [0:0] v_12343_0;
  wire [0:0] v_12344_0;
  reg [0:0] v_12345_0 = 1'h0;
  wire [0:0] v_12346_0;
  wire [0:0] v_12347_0;
  wire [0:0] _act_12348_0;
  wire [0:0] v_12349_0;
  wire [0:0] v_12350_0;
  wire [0:0] v_12351_0;
  wire [0:0] v_12352_0;
  wire [0:0] v_12353_0;
  wire [0:0] v_12354_0;
  reg [7:0] v_12356_0 = 8'h0;
  wire [7:0] v_12357_0;
  reg [7:0] v_12358_0 = 8'h0;
  wire [0:0] v_12359_0;
  wire [0:0] v_12360_0;
  wire [0:0] v_12361_0;
  wire [0:0] v_12362_0;
  wire [0:0] v_12363_0;
  wire [0:0] v_12364_0;
  wire [0:0] v_12365_0;
  wire [0:0] v_12366_0;
  wire [7:0] v_12367_0;
  wire [7:0] v_12368_0;
  wire [0:0] v_12369_0;
  wire [7:0] v_12370_0;
  wire [7:0] v_12371_0;
  wire [7:0] v_12372_0;
  wire [7:0] v_12373_0;
  // Instances
  //////////////////////////////////////////////////////////////////////////////
  assign v_1_0 = v_2_0 & v_6_0;
  assign v_2_0 = v_3_0 & v_12266_0;
  assign v_4_0 = v_5_0 & v_12265_0;
  assign v_5_0 = v_6_0 & v_95_0;
  assign v_6_0 = v_7_0 & v_30_0;
  assign v_7_0 = v_8_0 | v_12255_0;
  assign v_8_0 = 1'h1 & v_9_0;
  assign v_9_0 = v_10_0 == 16'h0;
  assign v_10_0 = v_11_0 ? v_12086_0 : v_12226_0;
  assign v_11_0 = 16'h1 < v_12_0;
  assign v_13_0 = v_14_0 & v_12083_0;
  assign v_14_0 = v_15_0 & v_34_0;
  assign v_15_0 = v_16_0 & v_12062_0;
  assign v_16_0 = 1'h1 & v_17_0;
  assign v_17_0 = ~v_18_0;
  assign v_19_0 = v_20_0 & v_12060_0;
  assign v_20_0 = ~v_21_0;
  assign v_21_0 = v_22_0 | v_689_0;
  assign v_22_0 = v_23_0 == 10'h0;
  assign v_24_0 = v_25_0 | v_587_0;
  assign v_25_0 = v_26_0 | v_4_0;
  assign v_26_0 = v_27_0 & v_30_0;
  assign v_27_0 = v_28_0 & 1'h1;
  assign v_28_0 = 1'h1 & v_29_0;
  assign v_29_0 = v_10_0 == 16'h0;
  assign v_30_0 = v_31_0 & v_586_0;
  assign v_31_0 = v_32_0 & v_33_0;
  assign v_32_0 = 1'h1 & v_18_0;
  assign v_33_0 = ~v_34_0;
  assign v_35_0 = v_36_0 | v_573_0;
  assign v_36_0 = v_37_0 | v_13_0;
  assign v_37_0 = v_38_0 & v_86_0;
  assign v_38_0 = v_39_0 & v_95_0;
  assign v_39_0 = v_40_0 & v_45_0;
  assign v_41_0 = v_13_0 | v_42_0;
  assign v_42_0 = v_43_0 | v_566_0;
  assign v_43_0 = v_44_0 & v_86_0;
  assign v_44_0 = ~v_45_0;
  assign v_45_0 = v_46_0 & v_564_0;
  assign v_46_0 = v_47_0 | v_321_0;
  assign v_47_0 = v_48_0 & v_320_0;
  assign v_48_0 = v_49_0 & 1'h1;
  assign v_49_0 = v_50_0 == 3'h7;
  assign v_50_0 = v_51_0 ? v_54_0 : v_271_0;
  assign v_51_0 = 16'h1 < v_52_0;
  assign v_53_0 = v_52_0 + 16'h1;
  assign v_55_0 = 1'h1 & v_56_0;
  assign v_56_0 = v_57_0 | v_177_0;
  assign v_57_0 = ~v_58_0;
  assign v_59_0 = v_60_0 | _act_63_0;
  assign v_61_0 = v_62_0 | v_173_0;
  assign v_62_0 = _act_63_0 & v_171_0;
  assign _act_63_0 = v_64_0 & 1'h1;
  assign v_64_0 = v_65_0 & v_66_0;
  assign v_65_0 = ~v_60_0;
  assign v_66_0 = ~v_67_0;
  assign v_68_0 = v_69_0 | v_166_0;
  assign v_69_0 = v_70_0 & v_163_0;
  assign v_70_0 = v_71_0 == v_78_0;
  assign v_71_0 = v_72_0 ? v_76_0 : v_77_0;
  assign v_72_0 = v_73_0 | v_74_0;
  assign v_73_0 = _act_63_0 ? 1'h1 : 1'h0;
  assign v_74_0 = v_75_0 ? 1'h0 : 1'h0;
  assign v_75_0 = ~_act_63_0;
  assign v_76_0 = v_77_0 + 5'h1;
  assign _act_79_0 = 1'h1 & _act_80_0;
  assign _act_80_0 = v_81_0 | v_136_0;
  assign v_81_0 = v_82_0 | v_127_0;
  assign v_82_0 = v_83_0 | v_125_0;
  assign v_83_0 = v_84_0 & v_51_0;
  assign v_84_0 = v_85_0 & v_121_0;
  assign v_85_0 = v_86_0 & v_115_0;
  assign v_86_0 = v_87_0 & v_91_0;
  assign v_87_0 = v_88_0 & v_90_0;
  assign v_88_0 = v_15_0 & v_89_0;
  assign v_89_0 = ~v_34_0;
  assign v_90_0 = ~v_34_0;
  assign v_92_0 = v_93_0 & v_95_0;
  assign v_93_0 = v_94_0 & v_87_0;
  assign v_94_0 = v_7_0 | v_91_0;
  assign v_95_0 = v_12_0 <= v_96_0;
  assign v_96_0 = v_97_0 + 16'h1;
  assign v_98_0 = v_99_0 | v_102_0;
  assign v_99_0 = v_100_0 | v_92_0;
  assign v_100_0 = v_93_0 & v_101_0;
  assign v_101_0 = ~v_95_0;
  assign v_102_0 = v_103_0 | v_4_0;
  assign v_103_0 = v_6_0 & v_104_0;
  assign v_104_0 = ~v_95_0;
  assign v_105_0 = v_106_0 | v_110_0;
  assign v_106_0 = v_107_0 | v_109_0;
  assign v_107_0 = v_100_0 ? v_108_0 : 16'h0;
  assign v_108_0 = v_97_0 + 16'h1;
  assign v_109_0 = v_92_0 ? 16'h0 : 16'h0;
  assign v_110_0 = v_111_0 | v_113_0;
  assign v_111_0 = v_103_0 ? v_112_0 : 16'h0;
  assign v_112_0 = v_97_0 + 16'h1;
  assign v_113_0 = v_4_0 ? 16'h0 : 16'h0;
  assign v_114_0 = ~v_91_0;
  assign v_115_0 = ~v_116_0;
  assign v_116_0 = v_117_0 | v_120_0;
  assign v_117_0 = v_118_0 & v_119_0;
  assign v_118_0 = v_46_0 & v_40_0;
  assign v_119_0 = v_10_0 == 16'h0;
  assign v_120_0 = v_121_0 & v_49_0;
  assign v_121_0 = v_122_0 & v_124_0;
  assign v_122_0 = v_123_0 & v_40_0;
  assign v_123_0 = ~v_46_0;
  assign v_124_0 = v_10_0 == 16'h0;
  assign v_125_0 = v_126_0 & v_51_0;
  assign v_126_0 = v_86_0 & v_116_0;
  assign v_127_0 = v_128_0 | v_129_0;
  assign v_128_0 = v_13_0 & v_51_0;
  assign v_129_0 = v_130_0 & v_51_0;
  assign v_130_0 = v_131_0 & v_135_0;
  assign v_131_0 = v_6_0 & v_132_0;
  assign v_132_0 = ~v_133_0;
  assign v_133_0 = 1'h0 | v_134_0;
  assign v_134_0 = 1'h0 & v_49_0;
  assign v_135_0 = ~1'h0;
  assign v_136_0 = v_137_0 | v_142_0;
  assign v_137_0 = v_138_0 | v_140_0;
  assign v_138_0 = v_139_0 & v_51_0;
  assign v_139_0 = v_131_0 & 1'h0;
  assign v_140_0 = v_141_0 & v_51_0;
  assign v_141_0 = v_6_0 & v_133_0;
  assign v_142_0 = v_143_0 | v_156_0;
  assign v_143_0 = v_144_0 | v_154_0;
  assign v_144_0 = v_145_0 & v_51_0;
  assign v_145_0 = v_146_0 & v_153_0;
  assign v_146_0 = v_147_0 & v_150_0;
  assign v_147_0 = v_94_0 & v_148_0;
  assign v_148_0 = v_87_0 & v_149_0;
  assign v_149_0 = ~v_91_0;
  assign v_150_0 = ~v_151_0;
  assign v_151_0 = 1'h0 | v_152_0;
  assign v_152_0 = 1'h0 & v_49_0;
  assign v_153_0 = ~1'h0;
  assign v_154_0 = v_155_0 & v_51_0;
  assign v_155_0 = v_146_0 & 1'h0;
  assign v_156_0 = v_157_0 | v_159_0;
  assign v_157_0 = v_158_0 & v_51_0;
  assign v_158_0 = v_147_0 & v_151_0;
  assign v_159_0 = v_160_0 & v_51_0;
  assign v_160_0 = v_85_0 & v_161_0;
  assign v_161_0 = ~v_121_0;
  assign v_162_0 = v_78_0 + 5'h1;
  assign v_163_0 = v_72_0 & v_164_0;
  assign v_164_0 = 1'h1 & v_165_0;
  assign v_165_0 = ~_act_80_0;
  assign v_166_0 = v_167_0 & _act_79_0;
  assign v_167_0 = ~v_72_0;
  assign v_168_0 = v_169_0 | v_170_0;
  assign v_169_0 = v_69_0 ? 1'h1 : 1'h0;
  assign v_170_0 = v_166_0 ? 1'h0 : 1'h0;
  assign v_171_0 = 1'h1 & v_172_0;
  assign v_172_0 = ~v_56_0;
  assign v_173_0 = v_60_0 & v_55_0;
  assign v_174_0 = v_175_0 | v_176_0;
  assign v_175_0 = v_62_0 ? 1'h1 : 1'h0;
  assign v_176_0 = v_173_0 ? _act_63_0 : 1'h0;
  assign v_177_0 = v_178_0 | v_183_0;
  assign v_178_0 = v_179_0 | v_181_0;
  assign v_179_0 = v_180_0 ? 1'h1 : 1'h0;
  assign v_180_0 = v_51_0 & v_147_0;
  assign v_181_0 = v_182_0 ? 1'h1 : 1'h0;
  assign v_182_0 = v_51_0 & v_86_0;
  assign v_183_0 = v_184_0 | v_186_0;
  assign v_184_0 = v_185_0 ? 1'h1 : 1'h0;
  assign v_185_0 = v_51_0 & v_6_0;
  assign v_186_0 = v_187_0 ? 1'h0 : 1'h0;
  assign v_187_0 = ~v_188_0;
  assign v_188_0 = v_185_0 | v_189_0;
  assign v_189_0 = v_180_0 | v_182_0;
  assign v_190_0 = v_60_0 ? v_191_0 : v_200_0;
  assign v_192_0 = v_193_0 & 1'h1;
  assign v_193_0 = v_194_0 | v_197_0;
  assign v_194_0 = v_195_0 ? 1'h0 : 1'h0;
  assign v_195_0 = ~v_196_0;
  assign v_196_0 = v_62_0 | v_173_0;
  assign v_197_0 = v_198_0 | v_199_0;
  assign v_198_0 = v_62_0 ? 1'h1 : 1'h0;
  assign v_199_0 = v_173_0 ? 1'h1 : 1'h0;
  assign v_200_0 = v_201_0 | v_269_0;
  assign v_201_0 = _act_63_0 ? v_202_0 : 3'h0;
  assign v_202_0 = v_203_0 ? v_218_0 : v_248_0;
  assign v_203_0 = v_204_0 & v_207_0;
  assign v_204_0 = v_205_0 & v_206_0;
  assign v_207_0 = v_208_0 == v_213_0;
  assign v_209_0 = v_210_0 | v_211_0;
  assign v_210_0 = 1'h1 ? v_71_0 : 5'h0;
  assign v_211_0 = v_212_0 ? 5'bxxxxx : 5'h0;
  assign v_212_0 = ~1'h1;
  assign v_214_0 = v_215_0 | v_216_0;
  assign v_215_0 = _act_79_0 ? v_78_0 : 5'h0;
  assign v_216_0 = v_217_0 ? 5'bxxxxx : 5'h0;
  assign v_217_0 = ~_act_79_0;
  assign v_219_0 = v_220_0 | v_246_0;
  assign v_220_0 = _act_79_0 ? v_221_0 : 3'h0;
  assign v_221_0 = v_222_0 | v_230_0;
  assign v_222_0 = v_223_0 | v_226_0;
  assign v_223_0 = v_224_0 | v_225_0;
  assign v_224_0 = v_128_0 ? 3'h0 : 3'h0;
  assign v_225_0 = v_129_0 ? v_50_0 : 3'h0;
  assign v_226_0 = v_227_0 | v_229_0;
  assign v_227_0 = v_138_0 ? v_228_0 : 3'h0;
  assign v_228_0 = v_50_0 + 3'h1;
  assign v_229_0 = v_140_0 ? 3'h0 : 3'h0;
  assign v_230_0 = v_231_0 | v_238_0;
  assign v_231_0 = v_232_0 | v_234_0;
  assign v_232_0 = v_233_0 ? 3'bxxx : 3'h0;
  assign v_233_0 = ~_act_80_0;
  assign v_234_0 = v_235_0 | v_236_0;
  assign v_235_0 = v_144_0 ? v_50_0 : 3'h0;
  assign v_236_0 = v_154_0 ? v_237_0 : 3'h0;
  assign v_237_0 = v_50_0 + 3'h1;
  assign v_238_0 = v_239_0 | v_242_0;
  assign v_239_0 = v_240_0 | v_241_0;
  assign v_240_0 = v_157_0 ? 3'h0 : 3'h0;
  assign v_241_0 = v_159_0 ? v_50_0 : 3'h0;
  assign v_242_0 = v_243_0 | v_245_0;
  assign v_243_0 = v_83_0 ? v_244_0 : 3'h0;
  assign v_244_0 = v_50_0 + 3'h1;
  assign v_245_0 = v_125_0 ? 3'h0 : 3'h0;
  assign v_246_0 = v_247_0 ? 3'bxxx : 3'h0;
  assign v_247_0 = ~_act_79_0;
  BlockRAMTrueDual#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(5), .DATA_WIDTH(3))
    ram248
      (.CLK(clock),
       .DI_A(v_253_0),
       .ADDR_A(v_249_0),
       .WE_A(v_255_0),
       .DO_A(v_248_0),
       .DI_B(v_261_0),
       .ADDR_B(v_257_0),
       .WE_B(v_265_0),
       .DO_B(v_248_1));
  assign v_249_0 = v_250_0 | v_251_0;
  assign v_250_0 = 1'h1 ? v_71_0 : 5'h0;
  assign v_251_0 = v_252_0 ? 5'bxxxxx : 5'h0;
  assign v_252_0 = ~1'h1;
  assign v_253_0 = v_254_0 ? 3'bxxx : 3'h0;
  assign v_254_0 = ~1'h0;
  assign v_255_0 = v_256_0 ? 1'h0 : 1'h0;
  assign v_256_0 = ~1'h0;
  assign v_257_0 = v_258_0 | v_259_0;
  assign v_258_0 = _act_79_0 ? v_78_0 : 5'h0;
  assign v_259_0 = v_260_0 ? 5'bxxxxx : 5'h0;
  assign v_260_0 = ~_act_79_0;
  assign v_261_0 = v_262_0 | v_263_0;
  assign v_262_0 = _act_79_0 ? v_221_0 : 3'h0;
  assign v_263_0 = v_264_0 ? 3'bxxx : 3'h0;
  assign v_264_0 = ~_act_79_0;
  assign v_265_0 = v_266_0 | v_267_0;
  assign v_266_0 = _act_79_0 ? 1'h1 : 1'h0;
  assign v_267_0 = v_268_0 ? 1'h0 : 1'h0;
  assign v_268_0 = ~_act_79_0;
  assign v_269_0 = v_270_0 ? 3'bxxx : 3'h0;
  assign v_270_0 = ~_act_63_0;
  assign v_272_0 = v_273_0 | v_284_0;
  assign v_273_0 = v_274_0 | v_279_0;
  assign v_274_0 = v_275_0 | v_277_0;
  assign v_275_0 = v_84_0 & v_276_0;
  assign v_276_0 = ~v_51_0;
  assign v_277_0 = v_126_0 & v_278_0;
  assign v_278_0 = ~v_51_0;
  assign v_279_0 = v_280_0 | v_282_0;
  assign v_280_0 = v_13_0 & v_281_0;
  assign v_281_0 = ~v_51_0;
  assign v_282_0 = v_130_0 & v_283_0;
  assign v_283_0 = ~v_51_0;
  assign v_284_0 = v_285_0 | v_290_0;
  assign v_285_0 = v_286_0 | v_288_0;
  assign v_286_0 = v_139_0 & v_287_0;
  assign v_287_0 = ~v_51_0;
  assign v_288_0 = v_141_0 & v_289_0;
  assign v_289_0 = ~v_51_0;
  assign v_290_0 = v_291_0 | v_296_0;
  assign v_291_0 = v_292_0 | v_294_0;
  assign v_292_0 = v_145_0 & v_293_0;
  assign v_293_0 = ~v_51_0;
  assign v_294_0 = v_155_0 & v_295_0;
  assign v_295_0 = ~v_51_0;
  assign v_296_0 = v_297_0 | v_299_0;
  assign v_297_0 = v_158_0 & v_298_0;
  assign v_298_0 = ~v_51_0;
  assign v_299_0 = v_160_0 & v_300_0;
  assign v_300_0 = ~v_51_0;
  assign v_301_0 = v_302_0 | v_309_0;
  assign v_302_0 = v_303_0 | v_306_0;
  assign v_303_0 = v_304_0 | v_305_0;
  assign v_304_0 = v_275_0 ? v_244_0 : 3'h0;
  assign v_305_0 = v_277_0 ? 3'h0 : 3'h0;
  assign v_306_0 = v_307_0 | v_308_0;
  assign v_307_0 = v_280_0 ? 3'h0 : 3'h0;
  assign v_308_0 = v_282_0 ? v_50_0 : 3'h0;
  assign v_309_0 = v_310_0 | v_313_0;
  assign v_310_0 = v_311_0 | v_312_0;
  assign v_311_0 = v_286_0 ? v_228_0 : 3'h0;
  assign v_312_0 = v_288_0 ? 3'h0 : 3'h0;
  assign v_313_0 = v_314_0 | v_317_0;
  assign v_314_0 = v_315_0 | v_316_0;
  assign v_315_0 = v_292_0 ? v_50_0 : 3'h0;
  assign v_316_0 = v_294_0 ? v_237_0 : 3'h0;
  assign v_317_0 = v_318_0 | v_319_0;
  assign v_318_0 = v_297_0 ? 3'h0 : 3'h0;
  assign v_319_0 = v_299_0 ? v_50_0 : 3'h0;
  assign v_320_0 = v_10_0 == 16'h0;
  assign v_321_0 = v_322_0 | v_324_0;
  assign v_322_0 = 1'h1 & v_323_0;
  assign v_323_0 = v_10_0 == 16'h1;
  assign v_324_0 = v_325_0 | 1'h0;
  assign v_325_0 = v_326_0 & v_563_0;
  assign v_326_0 = v_327_0 & 1'h1;
  assign v_327_0 = v_328_0 == 3'h7;
  assign v_328_0 = v_329_0 ? v_332_0 : v_514_0;
  assign v_329_0 = 16'h1 < v_330_0;
  assign v_331_0 = v_330_0 + 16'h1;
  assign v_333_0 = 1'h1 & v_334_0;
  assign v_334_0 = v_335_0 | v_420_0;
  assign v_335_0 = ~v_336_0;
  assign v_337_0 = v_338_0 | _act_341_0;
  assign v_339_0 = v_340_0 | v_416_0;
  assign v_340_0 = _act_341_0 & v_414_0;
  assign _act_341_0 = v_342_0 & 1'h1;
  assign v_342_0 = v_343_0 & v_344_0;
  assign v_343_0 = ~v_338_0;
  assign v_344_0 = ~v_345_0;
  assign v_346_0 = v_347_0 | v_409_0;
  assign v_347_0 = v_348_0 & v_406_0;
  assign v_348_0 = v_349_0 == v_356_0;
  assign v_349_0 = v_350_0 ? v_354_0 : v_355_0;
  assign v_350_0 = v_351_0 | v_352_0;
  assign v_351_0 = _act_341_0 ? 1'h1 : 1'h0;
  assign v_352_0 = v_353_0 ? 1'h0 : 1'h0;
  assign v_353_0 = ~_act_341_0;
  assign v_354_0 = v_355_0 + 5'h1;
  assign _act_357_0 = 1'h1 & _act_358_0;
  assign _act_358_0 = v_359_0 | v_382_0;
  assign v_359_0 = v_360_0 | v_373_0;
  assign v_360_0 = v_361_0 | v_371_0;
  assign v_361_0 = v_362_0 & v_329_0;
  assign v_362_0 = v_363_0 & v_369_0;
  assign v_363_0 = v_86_0 & v_364_0;
  assign v_364_0 = ~v_365_0;
  assign v_365_0 = v_366_0 | v_368_0;
  assign v_366_0 = v_118_0 & v_367_0;
  assign v_367_0 = v_10_0 == 16'h2;
  assign v_368_0 = v_369_0 & v_327_0;
  assign v_369_0 = v_122_0 & v_370_0;
  assign v_370_0 = v_10_0 == 16'h2;
  assign v_371_0 = v_372_0 & v_329_0;
  assign v_372_0 = v_86_0 & v_365_0;
  assign v_373_0 = v_374_0 | v_375_0;
  assign v_374_0 = v_13_0 & v_329_0;
  assign v_375_0 = v_376_0 & v_329_0;
  assign v_376_0 = v_377_0 & v_381_0;
  assign v_377_0 = v_6_0 & v_378_0;
  assign v_378_0 = ~v_379_0;
  assign v_379_0 = 1'h0 | v_380_0;
  assign v_380_0 = 1'h0 & v_327_0;
  assign v_381_0 = ~1'h0;
  assign v_382_0 = v_383_0 | v_388_0;
  assign v_383_0 = v_384_0 | v_386_0;
  assign v_384_0 = v_385_0 & v_329_0;
  assign v_385_0 = v_377_0 & 1'h0;
  assign v_386_0 = v_387_0 & v_329_0;
  assign v_387_0 = v_6_0 & v_379_0;
  assign v_388_0 = v_389_0 | v_399_0;
  assign v_389_0 = v_390_0 | v_397_0;
  assign v_390_0 = v_391_0 & v_329_0;
  assign v_391_0 = v_392_0 & v_396_0;
  assign v_392_0 = v_147_0 & v_393_0;
  assign v_393_0 = ~v_394_0;
  assign v_394_0 = 1'h0 | v_395_0;
  assign v_395_0 = 1'h0 & v_327_0;
  assign v_396_0 = ~1'h0;
  assign v_397_0 = v_398_0 & v_329_0;
  assign v_398_0 = v_392_0 & 1'h0;
  assign v_399_0 = v_400_0 | v_402_0;
  assign v_400_0 = v_401_0 & v_329_0;
  assign v_401_0 = v_147_0 & v_394_0;
  assign v_402_0 = v_403_0 & v_329_0;
  assign v_403_0 = v_363_0 & v_404_0;
  assign v_404_0 = ~v_369_0;
  assign v_405_0 = v_356_0 + 5'h1;
  assign v_406_0 = v_350_0 & v_407_0;
  assign v_407_0 = 1'h1 & v_408_0;
  assign v_408_0 = ~_act_358_0;
  assign v_409_0 = v_410_0 & _act_357_0;
  assign v_410_0 = ~v_350_0;
  assign v_411_0 = v_412_0 | v_413_0;
  assign v_412_0 = v_347_0 ? 1'h1 : 1'h0;
  assign v_413_0 = v_409_0 ? 1'h0 : 1'h0;
  assign v_414_0 = 1'h1 & v_415_0;
  assign v_415_0 = ~v_334_0;
  assign v_416_0 = v_338_0 & v_333_0;
  assign v_417_0 = v_418_0 | v_419_0;
  assign v_418_0 = v_340_0 ? 1'h1 : 1'h0;
  assign v_419_0 = v_416_0 ? _act_341_0 : 1'h0;
  assign v_420_0 = v_421_0 | v_426_0;
  assign v_421_0 = v_422_0 | v_424_0;
  assign v_422_0 = v_423_0 ? 1'h1 : 1'h0;
  assign v_423_0 = v_329_0 & v_147_0;
  assign v_424_0 = v_425_0 ? 1'h1 : 1'h0;
  assign v_425_0 = v_329_0 & v_86_0;
  assign v_426_0 = v_427_0 | v_429_0;
  assign v_427_0 = v_428_0 ? 1'h1 : 1'h0;
  assign v_428_0 = v_329_0 & v_6_0;
  assign v_429_0 = v_430_0 ? 1'h0 : 1'h0;
  assign v_430_0 = ~v_431_0;
  assign v_431_0 = v_428_0 | v_432_0;
  assign v_432_0 = v_423_0 | v_425_0;
  assign v_433_0 = v_338_0 ? v_434_0 : v_443_0;
  assign v_435_0 = v_436_0 & 1'h1;
  assign v_436_0 = v_437_0 | v_440_0;
  assign v_437_0 = v_438_0 ? 1'h0 : 1'h0;
  assign v_438_0 = ~v_439_0;
  assign v_439_0 = v_340_0 | v_416_0;
  assign v_440_0 = v_441_0 | v_442_0;
  assign v_441_0 = v_340_0 ? 1'h1 : 1'h0;
  assign v_442_0 = v_416_0 ? 1'h1 : 1'h0;
  assign v_443_0 = v_444_0 | v_512_0;
  assign v_444_0 = _act_341_0 ? v_445_0 : 3'h0;
  assign v_445_0 = v_446_0 ? v_461_0 : v_491_0;
  assign v_446_0 = v_447_0 & v_450_0;
  assign v_447_0 = v_448_0 & v_449_0;
  assign v_450_0 = v_451_0 == v_456_0;
  assign v_452_0 = v_453_0 | v_454_0;
  assign v_453_0 = 1'h1 ? v_349_0 : 5'h0;
  assign v_454_0 = v_455_0 ? 5'bxxxxx : 5'h0;
  assign v_455_0 = ~1'h1;
  assign v_457_0 = v_458_0 | v_459_0;
  assign v_458_0 = _act_357_0 ? v_356_0 : 5'h0;
  assign v_459_0 = v_460_0 ? 5'bxxxxx : 5'h0;
  assign v_460_0 = ~_act_357_0;
  assign v_462_0 = v_463_0 | v_489_0;
  assign v_463_0 = _act_357_0 ? v_464_0 : 3'h0;
  assign v_464_0 = v_465_0 | v_473_0;
  assign v_465_0 = v_466_0 | v_469_0;
  assign v_466_0 = v_467_0 | v_468_0;
  assign v_467_0 = v_374_0 ? 3'h0 : 3'h0;
  assign v_468_0 = v_375_0 ? v_328_0 : 3'h0;
  assign v_469_0 = v_470_0 | v_472_0;
  assign v_470_0 = v_384_0 ? v_471_0 : 3'h0;
  assign v_471_0 = v_328_0 + 3'h1;
  assign v_472_0 = v_386_0 ? 3'h0 : 3'h0;
  assign v_473_0 = v_474_0 | v_481_0;
  assign v_474_0 = v_475_0 | v_477_0;
  assign v_475_0 = v_476_0 ? 3'bxxx : 3'h0;
  assign v_476_0 = ~_act_358_0;
  assign v_477_0 = v_478_0 | v_479_0;
  assign v_478_0 = v_390_0 ? v_328_0 : 3'h0;
  assign v_479_0 = v_397_0 ? v_480_0 : 3'h0;
  assign v_480_0 = v_328_0 + 3'h1;
  assign v_481_0 = v_482_0 | v_485_0;
  assign v_482_0 = v_483_0 | v_484_0;
  assign v_483_0 = v_400_0 ? 3'h0 : 3'h0;
  assign v_484_0 = v_402_0 ? v_328_0 : 3'h0;
  assign v_485_0 = v_486_0 | v_488_0;
  assign v_486_0 = v_361_0 ? v_487_0 : 3'h0;
  assign v_487_0 = v_328_0 + 3'h1;
  assign v_488_0 = v_371_0 ? 3'h0 : 3'h0;
  assign v_489_0 = v_490_0 ? 3'bxxx : 3'h0;
  assign v_490_0 = ~_act_357_0;
  BlockRAMTrueDual#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(5), .DATA_WIDTH(3))
    ram491
      (.CLK(clock),
       .DI_A(v_496_0),
       .ADDR_A(v_492_0),
       .WE_A(v_498_0),
       .DO_A(v_491_0),
       .DI_B(v_504_0),
       .ADDR_B(v_500_0),
       .WE_B(v_508_0),
       .DO_B(v_491_1));
  assign v_492_0 = v_493_0 | v_494_0;
  assign v_493_0 = 1'h1 ? v_349_0 : 5'h0;
  assign v_494_0 = v_495_0 ? 5'bxxxxx : 5'h0;
  assign v_495_0 = ~1'h1;
  assign v_496_0 = v_497_0 ? 3'bxxx : 3'h0;
  assign v_497_0 = ~1'h0;
  assign v_498_0 = v_499_0 ? 1'h0 : 1'h0;
  assign v_499_0 = ~1'h0;
  assign v_500_0 = v_501_0 | v_502_0;
  assign v_501_0 = _act_357_0 ? v_356_0 : 5'h0;
  assign v_502_0 = v_503_0 ? 5'bxxxxx : 5'h0;
  assign v_503_0 = ~_act_357_0;
  assign v_504_0 = v_505_0 | v_506_0;
  assign v_505_0 = _act_357_0 ? v_464_0 : 3'h0;
  assign v_506_0 = v_507_0 ? 3'bxxx : 3'h0;
  assign v_507_0 = ~_act_357_0;
  assign v_508_0 = v_509_0 | v_510_0;
  assign v_509_0 = _act_357_0 ? 1'h1 : 1'h0;
  assign v_510_0 = v_511_0 ? 1'h0 : 1'h0;
  assign v_511_0 = ~_act_357_0;
  assign v_512_0 = v_513_0 ? 3'bxxx : 3'h0;
  assign v_513_0 = ~_act_341_0;
  assign v_515_0 = v_516_0 | v_527_0;
  assign v_516_0 = v_517_0 | v_522_0;
  assign v_517_0 = v_518_0 | v_520_0;
  assign v_518_0 = v_362_0 & v_519_0;
  assign v_519_0 = ~v_329_0;
  assign v_520_0 = v_372_0 & v_521_0;
  assign v_521_0 = ~v_329_0;
  assign v_522_0 = v_523_0 | v_525_0;
  assign v_523_0 = v_13_0 & v_524_0;
  assign v_524_0 = ~v_329_0;
  assign v_525_0 = v_376_0 & v_526_0;
  assign v_526_0 = ~v_329_0;
  assign v_527_0 = v_528_0 | v_533_0;
  assign v_528_0 = v_529_0 | v_531_0;
  assign v_529_0 = v_385_0 & v_530_0;
  assign v_530_0 = ~v_329_0;
  assign v_531_0 = v_387_0 & v_532_0;
  assign v_532_0 = ~v_329_0;
  assign v_533_0 = v_534_0 | v_539_0;
  assign v_534_0 = v_535_0 | v_537_0;
  assign v_535_0 = v_391_0 & v_536_0;
  assign v_536_0 = ~v_329_0;
  assign v_537_0 = v_398_0 & v_538_0;
  assign v_538_0 = ~v_329_0;
  assign v_539_0 = v_540_0 | v_542_0;
  assign v_540_0 = v_401_0 & v_541_0;
  assign v_541_0 = ~v_329_0;
  assign v_542_0 = v_403_0 & v_543_0;
  assign v_543_0 = ~v_329_0;
  assign v_544_0 = v_545_0 | v_552_0;
  assign v_545_0 = v_546_0 | v_549_0;
  assign v_546_0 = v_547_0 | v_548_0;
  assign v_547_0 = v_518_0 ? v_487_0 : 3'h0;
  assign v_548_0 = v_520_0 ? 3'h0 : 3'h0;
  assign v_549_0 = v_550_0 | v_551_0;
  assign v_550_0 = v_523_0 ? 3'h0 : 3'h0;
  assign v_551_0 = v_525_0 ? v_328_0 : 3'h0;
  assign v_552_0 = v_553_0 | v_556_0;
  assign v_553_0 = v_554_0 | v_555_0;
  assign v_554_0 = v_529_0 ? v_471_0 : 3'h0;
  assign v_555_0 = v_531_0 ? 3'h0 : 3'h0;
  assign v_556_0 = v_557_0 | v_560_0;
  assign v_557_0 = v_558_0 | v_559_0;
  assign v_558_0 = v_535_0 ? v_328_0 : 3'h0;
  assign v_559_0 = v_537_0 ? v_480_0 : 3'h0;
  assign v_560_0 = v_561_0 | v_562_0;
  assign v_561_0 = v_540_0 ? 3'h0 : 3'h0;
  assign v_562_0 = v_542_0 ? v_328_0 : 3'h0;
  assign v_563_0 = v_10_0 == 16'h2;
  assign v_564_0 = 16'h3 <= v_565_0;
  assign v_565_0 = v_10_0 + 16'h1;
  assign v_566_0 = v_92_0 & v_567_0;
  assign v_567_0 = ~v_91_0;
  assign v_568_0 = v_569_0 | v_570_0;
  assign v_569_0 = v_13_0 ? 1'h0 : 1'h0;
  assign v_570_0 = v_571_0 | v_572_0;
  assign v_571_0 = v_43_0 ? 1'h0 : 1'h0;
  assign v_572_0 = v_566_0 ? 1'h1 : 1'h0;
  assign v_573_0 = v_574_0 | v_575_0;
  assign v_574_0 = v_5_0 & v_3_0;
  assign v_575_0 = v_31_0 & v_576_0;
  assign v_576_0 = v_577_0 & v_3_0;
  assign v_577_0 = v_578_0 < v_97_0;
  assign v_579_0 = v_580_0 | v_583_0;
  assign v_580_0 = v_581_0 | v_582_0;
  assign v_581_0 = v_37_0 ? 1'h1 : 1'h0;
  assign v_582_0 = v_13_0 ? 1'h0 : 1'h0;
  assign v_583_0 = v_584_0 | v_585_0;
  assign v_584_0 = v_574_0 ? 1'h1 : 1'h0;
  assign v_585_0 = v_575_0 ? 1'h1 : 1'h0;
  assign v_586_0 = ~v_576_0;
  assign v_587_0 = v_588_0 | v_675_0;
  assign v_588_0 = v_589_0 | v_601_0;
  assign v_589_0 = v_590_0 & v_148_0;
  assign v_590_0 = v_591_0 & v_593_0;
  assign v_591_0 = 1'h1 & v_592_0;
  assign v_592_0 = v_10_0 == 16'h1;
  assign v_593_0 = v_594_0 & v_595_0;
  assign v_594_0 = ~v_22_0;
  assign v_595_0 = ~v_596_0;
  assign v_596_0 = v_597_0 == 10'h0;
  assign v_598_0 = v_599_0 | v_611_0;
  assign v_599_0 = v_600_0 | v_605_0;
  assign v_600_0 = v_589_0 | v_601_0;
  assign v_601_0 = v_602_0 & v_148_0;
  assign v_602_0 = v_603_0 & 1'h1;
  assign v_603_0 = 1'h1 & v_604_0;
  assign v_604_0 = v_10_0 == 16'h0;
  assign v_605_0 = v_606_0 | v_607_0;
  assign v_606_0 = v_92_0 & v_91_0;
  assign v_607_0 = v_608_0 & v_30_0;
  assign v_608_0 = v_609_0 & v_593_0;
  assign v_609_0 = 1'h1 & v_610_0;
  assign v_610_0 = v_10_0 == 16'h1;
  assign v_611_0 = v_612_0 | v_613_0;
  assign v_612_0 = v_26_0 | v_4_0;
  assign v_613_0 = v_614_0 | v_656_0;
  assign v_614_0 = v_615_0 & 1'h1;
  assign v_617_0 = v_618_0 | v_648_0;
  assign v_618_0 = v_619_0 | v_623_0;
  assign v_619_0 = v_620_0 & v_148_0;
  assign v_621_0 = v_622_0 | v_630_0;
  assign v_622_0 = v_619_0 | v_623_0;
  assign v_623_0 = v_624_0 & v_148_0;
  assign v_624_0 = v_625_0 & v_629_0;
  assign v_625_0 = v_626_0 & v_628_0;
  assign v_626_0 = 1'h1 & v_627_0;
  assign v_627_0 = v_10_0 == 16'h2;
  assign v_628_0 = ~v_596_0;
  assign v_629_0 = ~v_620_0;
  assign v_630_0 = v_631_0 | v_632_0;
  assign v_631_0 = v_620_0 & v_30_0;
  assign v_632_0 = v_633_0 & v_30_0;
  assign v_633_0 = v_634_0 & v_637_0;
  assign v_634_0 = v_635_0 & v_628_0;
  assign v_635_0 = 1'h1 & v_636_0;
  assign v_636_0 = v_10_0 == 16'h2;
  assign v_637_0 = ~v_620_0;
  assign v_638_0 = v_639_0 | v_644_0;
  assign v_639_0 = v_640_0 | v_643_0;
  assign v_640_0 = v_619_0 ? v_641_0 : 1'h0;
  assign v_641_0 = ~v_642_0;
  assign v_643_0 = v_623_0 ? 1'h1 : 1'h0;
  assign v_644_0 = v_645_0 | v_647_0;
  assign v_645_0 = v_631_0 ? v_646_0 : 1'h0;
  assign v_646_0 = ~v_642_0;
  assign v_647_0 = v_632_0 ? 1'h1 : 1'h0;
  assign v_648_0 = v_631_0 | v_632_0;
  assign v_649_0 = v_650_0 | v_653_0;
  assign v_650_0 = v_651_0 | v_652_0;
  assign v_651_0 = v_619_0 ? 1'h0 : 1'h0;
  assign v_652_0 = v_623_0 ? 1'h1 : 1'h0;
  assign v_653_0 = v_654_0 | v_655_0;
  assign v_654_0 = v_631_0 ? 1'h0 : 1'h0;
  assign v_655_0 = v_632_0 ? 1'h1 : 1'h0;
  assign v_656_0 = v_616_0 & 1'h1;
  assign v_657_0 = v_658_0 | v_667_0;
  assign v_658_0 = v_659_0 | v_664_0;
  assign v_659_0 = v_660_0 | v_662_0;
  assign v_660_0 = v_589_0 ? v_661_0 : 10'h0;
  assign v_661_0 = v_597_0 - 10'h1;
  assign v_662_0 = v_601_0 ? v_663_0 : 10'h0;
  assign v_663_0 = v_597_0 + 10'h1;
  assign v_664_0 = v_665_0 | v_666_0;
  assign v_665_0 = v_606_0 ? 10'h0 : 10'h0;
  assign v_666_0 = v_607_0 ? v_661_0 : 10'h0;
  assign v_667_0 = v_668_0 | v_671_0;
  assign v_668_0 = v_669_0 | v_670_0;
  assign v_669_0 = v_26_0 ? v_663_0 : 10'h0;
  assign v_670_0 = v_4_0 ? 10'h0 : 10'h0;
  assign v_671_0 = v_672_0 | v_673_0;
  assign v_672_0 = v_614_0 ? v_661_0 : 10'h0;
  assign v_673_0 = v_656_0 ? v_674_0 : 10'h0;
  assign v_674_0 = v_597_0 + 10'h1;
  assign v_675_0 = v_606_0 | v_607_0;
  assign v_676_0 = v_677_0 | v_681_0;
  assign v_677_0 = v_678_0 | v_680_0;
  assign v_678_0 = v_26_0 ? v_679_0 : 10'h0;
  assign v_679_0 = v_23_0 + 10'h1;
  assign v_680_0 = v_4_0 ? 10'h0 : 10'h0;
  assign v_681_0 = v_682_0 | v_686_0;
  assign v_682_0 = v_683_0 | v_685_0;
  assign v_683_0 = v_589_0 ? v_684_0 : 10'h0;
  assign v_684_0 = v_23_0 - 10'h1;
  assign v_685_0 = v_601_0 ? v_679_0 : 10'h0;
  assign v_686_0 = v_687_0 | v_688_0;
  assign v_687_0 = v_606_0 ? 10'h0 : 10'h0;
  assign v_688_0 = v_607_0 ? v_684_0 : 10'h0;
  assign v_689_0 = v_690_0 == v_11948_0;
  assign v_691_0 = v_692_0 | v_693_0;
  assign v_692_0 = v_589_0 | v_601_0;
  assign v_693_0 = v_607_0 | v_26_0;
  assign v_694_0 = v_695_0 | v_11945_0;
  assign v_695_0 = v_696_0 | v_11944_0;
  assign v_696_0 = v_589_0 ? v_697_0 : 3'h0;
  assign v_698_0 = v_699_0 | v_700_0;
  assign v_699_0 = v_589_0 | v_601_0;
  assign v_700_0 = v_607_0 | v_26_0;
  assign v_701_0 = v_702_0 | v_11941_0;
  assign v_702_0 = v_703_0 | v_11940_0;
  assign v_703_0 = v_589_0 ? v_704_0 : 3'h0;
  assign v_705_0 = v_706_0 | v_707_0;
  assign v_706_0 = v_589_0 | v_601_0;
  assign v_707_0 = v_607_0 | v_26_0;
  assign v_708_0 = v_709_0 | v_11937_0;
  assign v_709_0 = v_710_0 | v_11936_0;
  assign v_710_0 = v_589_0 ? v_711_0 : 3'h0;
  assign v_712_0 = v_713_0 | v_714_0;
  assign v_713_0 = v_589_0 | v_601_0;
  assign v_714_0 = v_607_0 | v_26_0;
  assign v_715_0 = v_716_0 | v_11933_0;
  assign v_716_0 = v_717_0 | v_11932_0;
  assign v_717_0 = v_589_0 ? v_718_0 : 3'h0;
  assign v_719_0 = v_720_0 | v_721_0;
  assign v_720_0 = v_589_0 | v_601_0;
  assign v_721_0 = v_607_0 | v_26_0;
  assign v_722_0 = v_723_0 | v_11929_0;
  assign v_723_0 = v_724_0 | v_11928_0;
  assign v_724_0 = v_589_0 ? v_725_0 : 3'h0;
  assign v_726_0 = v_727_0 | v_728_0;
  assign v_727_0 = v_589_0 | v_601_0;
  assign v_728_0 = v_607_0 | v_26_0;
  assign v_729_0 = v_730_0 | v_11925_0;
  assign v_730_0 = v_731_0 | v_11924_0;
  assign v_731_0 = v_589_0 ? v_732_0 : 3'h0;
  assign v_733_0 = v_734_0 | v_735_0;
  assign v_734_0 = v_589_0 | v_601_0;
  assign v_735_0 = v_607_0 | v_26_0;
  assign v_736_0 = v_737_0 | v_11921_0;
  assign v_737_0 = v_738_0 | v_11920_0;
  assign v_738_0 = v_589_0 ? v_739_0 : 3'h0;
  assign v_740_0 = v_741_0 | v_742_0;
  assign v_741_0 = v_589_0 | v_601_0;
  assign v_742_0 = v_607_0 | v_26_0;
  assign v_743_0 = v_744_0 | v_11917_0;
  assign v_744_0 = v_745_0 | v_11916_0;
  assign v_745_0 = v_589_0 ? v_746_0 : 3'h0;
  assign v_747_0 = v_748_0 | v_749_0;
  assign v_748_0 = v_589_0 | v_601_0;
  assign v_749_0 = v_607_0 | v_26_0;
  assign v_750_0 = v_751_0 | v_11913_0;
  assign v_751_0 = v_752_0 | v_11912_0;
  assign v_752_0 = v_589_0 ? v_753_0 : 3'h0;
  assign v_754_0 = v_755_0 | v_756_0;
  assign v_755_0 = v_589_0 | v_601_0;
  assign v_756_0 = v_607_0 | v_26_0;
  assign v_757_0 = v_758_0 | v_11909_0;
  assign v_758_0 = v_759_0 | v_11908_0;
  assign v_759_0 = v_589_0 ? v_760_0 : 3'h0;
  assign v_761_0 = v_762_0 | v_763_0;
  assign v_762_0 = v_589_0 | v_601_0;
  assign v_763_0 = v_607_0 | v_26_0;
  assign v_764_0 = v_765_0 | v_11905_0;
  assign v_765_0 = v_766_0 | v_11904_0;
  assign v_766_0 = v_589_0 ? v_767_0 : 3'h0;
  assign v_768_0 = v_769_0 | v_770_0;
  assign v_769_0 = v_589_0 | v_601_0;
  assign v_770_0 = v_607_0 | v_26_0;
  assign v_771_0 = v_772_0 | v_11901_0;
  assign v_772_0 = v_773_0 | v_11900_0;
  assign v_773_0 = v_589_0 ? v_774_0 : 3'h0;
  assign v_775_0 = v_776_0 | v_777_0;
  assign v_776_0 = v_589_0 | v_601_0;
  assign v_777_0 = v_607_0 | v_26_0;
  assign v_778_0 = v_779_0 | v_11897_0;
  assign v_779_0 = v_780_0 | v_11896_0;
  assign v_780_0 = v_589_0 ? v_781_0 : 3'h0;
  assign v_782_0 = v_783_0 | v_784_0;
  assign v_783_0 = v_589_0 | v_601_0;
  assign v_784_0 = v_607_0 | v_26_0;
  assign v_785_0 = v_786_0 | v_11893_0;
  assign v_786_0 = v_787_0 | v_11892_0;
  assign v_787_0 = v_589_0 ? v_788_0 : 3'h0;
  assign v_789_0 = v_790_0 | v_791_0;
  assign v_790_0 = v_589_0 | v_601_0;
  assign v_791_0 = v_607_0 | v_26_0;
  assign v_792_0 = v_793_0 | v_11889_0;
  assign v_793_0 = v_794_0 | v_11888_0;
  assign v_794_0 = v_589_0 ? v_795_0 : 3'h0;
  assign v_796_0 = v_797_0 | v_798_0;
  assign v_797_0 = v_589_0 | v_601_0;
  assign v_798_0 = v_607_0 | v_26_0;
  assign v_799_0 = v_800_0 | v_11885_0;
  assign v_800_0 = v_801_0 | v_11884_0;
  assign v_801_0 = v_589_0 ? v_802_0 : 3'h0;
  assign v_803_0 = v_804_0 | v_805_0;
  assign v_804_0 = v_589_0 | v_601_0;
  assign v_805_0 = v_607_0 | v_26_0;
  assign v_806_0 = v_807_0 | v_11881_0;
  assign v_807_0 = v_808_0 | v_11880_0;
  assign v_808_0 = v_589_0 ? v_809_0 : 3'h0;
  assign v_810_0 = v_811_0 | v_812_0;
  assign v_811_0 = v_589_0 | v_601_0;
  assign v_812_0 = v_607_0 | v_26_0;
  assign v_813_0 = v_814_0 | v_11877_0;
  assign v_814_0 = v_815_0 | v_11876_0;
  assign v_815_0 = v_589_0 ? v_816_0 : 3'h0;
  assign v_817_0 = v_818_0 | v_819_0;
  assign v_818_0 = v_589_0 | v_601_0;
  assign v_819_0 = v_607_0 | v_26_0;
  assign v_820_0 = v_821_0 | v_11873_0;
  assign v_821_0 = v_822_0 | v_11872_0;
  assign v_822_0 = v_589_0 ? v_823_0 : 3'h0;
  assign v_824_0 = v_825_0 | v_826_0;
  assign v_825_0 = v_589_0 | v_601_0;
  assign v_826_0 = v_607_0 | v_26_0;
  assign v_827_0 = v_828_0 | v_11869_0;
  assign v_828_0 = v_829_0 | v_11868_0;
  assign v_829_0 = v_589_0 ? v_830_0 : 3'h0;
  assign v_831_0 = v_832_0 | v_833_0;
  assign v_832_0 = v_589_0 | v_601_0;
  assign v_833_0 = v_607_0 | v_26_0;
  assign v_834_0 = v_835_0 | v_11865_0;
  assign v_835_0 = v_836_0 | v_11864_0;
  assign v_836_0 = v_589_0 ? v_837_0 : 3'h0;
  assign v_838_0 = v_839_0 | v_840_0;
  assign v_839_0 = v_589_0 | v_601_0;
  assign v_840_0 = v_607_0 | v_26_0;
  assign v_841_0 = v_842_0 | v_11861_0;
  assign v_842_0 = v_843_0 | v_11860_0;
  assign v_843_0 = v_589_0 ? v_844_0 : 3'h0;
  assign v_845_0 = v_846_0 | v_847_0;
  assign v_846_0 = v_589_0 | v_601_0;
  assign v_847_0 = v_607_0 | v_26_0;
  assign v_848_0 = v_849_0 | v_11857_0;
  assign v_849_0 = v_850_0 | v_11856_0;
  assign v_850_0 = v_589_0 ? v_851_0 : 3'h0;
  assign v_852_0 = v_853_0 | v_854_0;
  assign v_853_0 = v_589_0 | v_601_0;
  assign v_854_0 = v_607_0 | v_26_0;
  assign v_855_0 = v_856_0 | v_11853_0;
  assign v_856_0 = v_857_0 | v_11852_0;
  assign v_857_0 = v_589_0 ? v_858_0 : 3'h0;
  assign v_859_0 = v_860_0 | v_861_0;
  assign v_860_0 = v_589_0 | v_601_0;
  assign v_861_0 = v_607_0 | v_26_0;
  assign v_862_0 = v_863_0 | v_11849_0;
  assign v_863_0 = v_864_0 | v_11848_0;
  assign v_864_0 = v_589_0 ? v_865_0 : 3'h0;
  assign v_866_0 = v_867_0 | v_868_0;
  assign v_867_0 = v_589_0 | v_601_0;
  assign v_868_0 = v_607_0 | v_26_0;
  assign v_869_0 = v_870_0 | v_11845_0;
  assign v_870_0 = v_871_0 | v_11844_0;
  assign v_871_0 = v_589_0 ? v_872_0 : 3'h0;
  assign v_873_0 = v_874_0 | v_875_0;
  assign v_874_0 = v_589_0 | v_601_0;
  assign v_875_0 = v_607_0 | v_26_0;
  assign v_876_0 = v_877_0 | v_11841_0;
  assign v_877_0 = v_878_0 | v_11840_0;
  assign v_878_0 = v_589_0 ? v_879_0 : 3'h0;
  assign v_880_0 = v_881_0 | v_882_0;
  assign v_881_0 = v_589_0 | v_601_0;
  assign v_882_0 = v_607_0 | v_26_0;
  assign v_883_0 = v_884_0 | v_11837_0;
  assign v_884_0 = v_885_0 | v_11836_0;
  assign v_885_0 = v_589_0 ? v_886_0 : 3'h0;
  assign v_887_0 = v_888_0 | v_889_0;
  assign v_888_0 = v_589_0 | v_601_0;
  assign v_889_0 = v_607_0 | v_26_0;
  assign v_890_0 = v_891_0 | v_11833_0;
  assign v_891_0 = v_892_0 | v_11832_0;
  assign v_892_0 = v_589_0 ? v_893_0 : 3'h0;
  assign v_894_0 = v_895_0 | v_896_0;
  assign v_895_0 = v_589_0 | v_601_0;
  assign v_896_0 = v_607_0 | v_26_0;
  assign v_897_0 = v_898_0 | v_11829_0;
  assign v_898_0 = v_899_0 | v_11828_0;
  assign v_899_0 = v_589_0 ? v_900_0 : 3'h0;
  assign v_901_0 = v_902_0 | v_903_0;
  assign v_902_0 = v_589_0 | v_601_0;
  assign v_903_0 = v_607_0 | v_26_0;
  assign v_904_0 = v_905_0 | v_11825_0;
  assign v_905_0 = v_906_0 | v_11824_0;
  assign v_906_0 = v_589_0 ? v_907_0 : 3'h0;
  assign v_908_0 = v_909_0 | v_910_0;
  assign v_909_0 = v_589_0 | v_601_0;
  assign v_910_0 = v_607_0 | v_26_0;
  assign v_911_0 = v_912_0 | v_11821_0;
  assign v_912_0 = v_913_0 | v_11820_0;
  assign v_913_0 = v_589_0 ? v_914_0 : 3'h0;
  assign v_915_0 = v_916_0 | v_917_0;
  assign v_916_0 = v_589_0 | v_601_0;
  assign v_917_0 = v_607_0 | v_26_0;
  assign v_918_0 = v_919_0 | v_11817_0;
  assign v_919_0 = v_920_0 | v_11816_0;
  assign v_920_0 = v_589_0 ? v_921_0 : 3'h0;
  assign v_922_0 = v_923_0 | v_924_0;
  assign v_923_0 = v_589_0 | v_601_0;
  assign v_924_0 = v_607_0 | v_26_0;
  assign v_925_0 = v_926_0 | v_11813_0;
  assign v_926_0 = v_927_0 | v_11812_0;
  assign v_927_0 = v_589_0 ? v_928_0 : 3'h0;
  assign v_929_0 = v_930_0 | v_931_0;
  assign v_930_0 = v_589_0 | v_601_0;
  assign v_931_0 = v_607_0 | v_26_0;
  assign v_932_0 = v_933_0 | v_11809_0;
  assign v_933_0 = v_934_0 | v_11808_0;
  assign v_934_0 = v_589_0 ? v_935_0 : 3'h0;
  assign v_936_0 = v_937_0 | v_938_0;
  assign v_937_0 = v_589_0 | v_601_0;
  assign v_938_0 = v_607_0 | v_26_0;
  assign v_939_0 = v_940_0 | v_11805_0;
  assign v_940_0 = v_941_0 | v_11804_0;
  assign v_941_0 = v_589_0 ? v_942_0 : 3'h0;
  assign v_943_0 = v_944_0 | v_945_0;
  assign v_944_0 = v_589_0 | v_601_0;
  assign v_945_0 = v_607_0 | v_26_0;
  assign v_946_0 = v_947_0 | v_11801_0;
  assign v_947_0 = v_948_0 | v_11800_0;
  assign v_948_0 = v_589_0 ? v_949_0 : 3'h0;
  assign v_950_0 = v_951_0 | v_952_0;
  assign v_951_0 = v_589_0 | v_601_0;
  assign v_952_0 = v_607_0 | v_26_0;
  assign v_953_0 = v_954_0 | v_11797_0;
  assign v_954_0 = v_955_0 | v_11796_0;
  assign v_955_0 = v_589_0 ? v_956_0 : 3'h0;
  assign v_957_0 = v_958_0 | v_959_0;
  assign v_958_0 = v_589_0 | v_601_0;
  assign v_959_0 = v_607_0 | v_26_0;
  assign v_960_0 = v_961_0 | v_11793_0;
  assign v_961_0 = v_962_0 | v_11792_0;
  assign v_962_0 = v_589_0 ? v_963_0 : 3'h0;
  assign v_964_0 = v_965_0 | v_966_0;
  assign v_965_0 = v_589_0 | v_601_0;
  assign v_966_0 = v_607_0 | v_26_0;
  assign v_967_0 = v_968_0 | v_11789_0;
  assign v_968_0 = v_969_0 | v_11788_0;
  assign v_969_0 = v_589_0 ? v_970_0 : 3'h0;
  assign v_971_0 = v_972_0 | v_973_0;
  assign v_972_0 = v_589_0 | v_601_0;
  assign v_973_0 = v_607_0 | v_26_0;
  assign v_974_0 = v_975_0 | v_11785_0;
  assign v_975_0 = v_976_0 | v_11784_0;
  assign v_976_0 = v_589_0 ? v_977_0 : 3'h0;
  assign v_978_0 = v_979_0 | v_980_0;
  assign v_979_0 = v_589_0 | v_601_0;
  assign v_980_0 = v_607_0 | v_26_0;
  assign v_981_0 = v_982_0 | v_11781_0;
  assign v_982_0 = v_983_0 | v_11780_0;
  assign v_983_0 = v_589_0 ? v_984_0 : 3'h0;
  assign v_985_0 = v_986_0 | v_987_0;
  assign v_986_0 = v_589_0 | v_601_0;
  assign v_987_0 = v_607_0 | v_26_0;
  assign v_988_0 = v_989_0 | v_11777_0;
  assign v_989_0 = v_990_0 | v_11776_0;
  assign v_990_0 = v_589_0 ? v_991_0 : 3'h0;
  assign v_992_0 = v_993_0 | v_994_0;
  assign v_993_0 = v_589_0 | v_601_0;
  assign v_994_0 = v_607_0 | v_26_0;
  assign v_995_0 = v_996_0 | v_11773_0;
  assign v_996_0 = v_997_0 | v_11772_0;
  assign v_997_0 = v_589_0 ? v_998_0 : 3'h0;
  assign v_999_0 = v_1000_0 | v_1001_0;
  assign v_1000_0 = v_589_0 | v_601_0;
  assign v_1001_0 = v_607_0 | v_26_0;
  assign v_1002_0 = v_1003_0 | v_11769_0;
  assign v_1003_0 = v_1004_0 | v_11768_0;
  assign v_1004_0 = v_589_0 ? v_1005_0 : 3'h0;
  assign v_1006_0 = v_1007_0 | v_1008_0;
  assign v_1007_0 = v_589_0 | v_601_0;
  assign v_1008_0 = v_607_0 | v_26_0;
  assign v_1009_0 = v_1010_0 | v_11765_0;
  assign v_1010_0 = v_1011_0 | v_11764_0;
  assign v_1011_0 = v_589_0 ? v_1012_0 : 3'h0;
  assign v_1013_0 = v_1014_0 | v_1015_0;
  assign v_1014_0 = v_589_0 | v_601_0;
  assign v_1015_0 = v_607_0 | v_26_0;
  assign v_1016_0 = v_1017_0 | v_11761_0;
  assign v_1017_0 = v_1018_0 | v_11760_0;
  assign v_1018_0 = v_589_0 ? v_1019_0 : 3'h0;
  assign v_1020_0 = v_1021_0 | v_1022_0;
  assign v_1021_0 = v_589_0 | v_601_0;
  assign v_1022_0 = v_607_0 | v_26_0;
  assign v_1023_0 = v_1024_0 | v_11757_0;
  assign v_1024_0 = v_1025_0 | v_11756_0;
  assign v_1025_0 = v_589_0 ? v_1026_0 : 3'h0;
  assign v_1027_0 = v_1028_0 | v_1029_0;
  assign v_1028_0 = v_589_0 | v_601_0;
  assign v_1029_0 = v_607_0 | v_26_0;
  assign v_1030_0 = v_1031_0 | v_11753_0;
  assign v_1031_0 = v_1032_0 | v_11752_0;
  assign v_1032_0 = v_589_0 ? v_1033_0 : 3'h0;
  assign v_1034_0 = v_1035_0 | v_1036_0;
  assign v_1035_0 = v_589_0 | v_601_0;
  assign v_1036_0 = v_607_0 | v_26_0;
  assign v_1037_0 = v_1038_0 | v_11749_0;
  assign v_1038_0 = v_1039_0 | v_11748_0;
  assign v_1039_0 = v_589_0 ? v_1040_0 : 3'h0;
  assign v_1041_0 = v_1042_0 | v_1043_0;
  assign v_1042_0 = v_589_0 | v_601_0;
  assign v_1043_0 = v_607_0 | v_26_0;
  assign v_1044_0 = v_1045_0 | v_11745_0;
  assign v_1045_0 = v_1046_0 | v_11744_0;
  assign v_1046_0 = v_589_0 ? v_1047_0 : 3'h0;
  assign v_1048_0 = v_1049_0 | v_1050_0;
  assign v_1049_0 = v_589_0 | v_601_0;
  assign v_1050_0 = v_607_0 | v_26_0;
  assign v_1051_0 = v_1052_0 | v_11741_0;
  assign v_1052_0 = v_1053_0 | v_11740_0;
  assign v_1053_0 = v_589_0 ? v_1054_0 : 3'h0;
  assign v_1055_0 = v_1056_0 | v_1057_0;
  assign v_1056_0 = v_589_0 | v_601_0;
  assign v_1057_0 = v_607_0 | v_26_0;
  assign v_1058_0 = v_1059_0 | v_11737_0;
  assign v_1059_0 = v_1060_0 | v_11736_0;
  assign v_1060_0 = v_589_0 ? v_1061_0 : 3'h0;
  assign v_1062_0 = v_1063_0 | v_1064_0;
  assign v_1063_0 = v_589_0 | v_601_0;
  assign v_1064_0 = v_607_0 | v_26_0;
  assign v_1065_0 = v_1066_0 | v_11733_0;
  assign v_1066_0 = v_1067_0 | v_11732_0;
  assign v_1067_0 = v_589_0 ? v_1068_0 : 3'h0;
  assign v_1069_0 = v_1070_0 | v_1071_0;
  assign v_1070_0 = v_589_0 | v_601_0;
  assign v_1071_0 = v_607_0 | v_26_0;
  assign v_1072_0 = v_1073_0 | v_11729_0;
  assign v_1073_0 = v_1074_0 | v_11728_0;
  assign v_1074_0 = v_589_0 ? v_1075_0 : 3'h0;
  assign v_1076_0 = v_1077_0 | v_1078_0;
  assign v_1077_0 = v_589_0 | v_601_0;
  assign v_1078_0 = v_607_0 | v_26_0;
  assign v_1079_0 = v_1080_0 | v_11725_0;
  assign v_1080_0 = v_1081_0 | v_11724_0;
  assign v_1081_0 = v_589_0 ? v_1082_0 : 3'h0;
  assign v_1083_0 = v_1084_0 | v_1085_0;
  assign v_1084_0 = v_589_0 | v_601_0;
  assign v_1085_0 = v_607_0 | v_26_0;
  assign v_1086_0 = v_1087_0 | v_11721_0;
  assign v_1087_0 = v_1088_0 | v_11720_0;
  assign v_1088_0 = v_589_0 ? v_1089_0 : 3'h0;
  assign v_1090_0 = v_1091_0 | v_1092_0;
  assign v_1091_0 = v_589_0 | v_601_0;
  assign v_1092_0 = v_607_0 | v_26_0;
  assign v_1093_0 = v_1094_0 | v_11717_0;
  assign v_1094_0 = v_1095_0 | v_11716_0;
  assign v_1095_0 = v_589_0 ? v_1096_0 : 3'h0;
  assign v_1097_0 = v_1098_0 | v_1099_0;
  assign v_1098_0 = v_589_0 | v_601_0;
  assign v_1099_0 = v_607_0 | v_26_0;
  assign v_1100_0 = v_1101_0 | v_11713_0;
  assign v_1101_0 = v_1102_0 | v_11712_0;
  assign v_1102_0 = v_589_0 ? v_1103_0 : 3'h0;
  assign v_1104_0 = v_1105_0 | v_1106_0;
  assign v_1105_0 = v_589_0 | v_601_0;
  assign v_1106_0 = v_607_0 | v_26_0;
  assign v_1107_0 = v_1108_0 | v_11709_0;
  assign v_1108_0 = v_1109_0 | v_11708_0;
  assign v_1109_0 = v_589_0 ? v_1110_0 : 3'h0;
  assign v_1111_0 = v_1112_0 | v_1113_0;
  assign v_1112_0 = v_589_0 | v_601_0;
  assign v_1113_0 = v_607_0 | v_26_0;
  assign v_1114_0 = v_1115_0 | v_11705_0;
  assign v_1115_0 = v_1116_0 | v_11704_0;
  assign v_1116_0 = v_589_0 ? v_1117_0 : 3'h0;
  assign v_1118_0 = v_1119_0 | v_1120_0;
  assign v_1119_0 = v_589_0 | v_601_0;
  assign v_1120_0 = v_607_0 | v_26_0;
  assign v_1121_0 = v_1122_0 | v_11701_0;
  assign v_1122_0 = v_1123_0 | v_11700_0;
  assign v_1123_0 = v_589_0 ? v_1124_0 : 3'h0;
  assign v_1125_0 = v_1126_0 | v_1127_0;
  assign v_1126_0 = v_589_0 | v_601_0;
  assign v_1127_0 = v_607_0 | v_26_0;
  assign v_1128_0 = v_1129_0 | v_11697_0;
  assign v_1129_0 = v_1130_0 | v_11696_0;
  assign v_1130_0 = v_589_0 ? v_1131_0 : 3'h0;
  assign v_1132_0 = v_1133_0 | v_1134_0;
  assign v_1133_0 = v_589_0 | v_601_0;
  assign v_1134_0 = v_607_0 | v_26_0;
  assign v_1135_0 = v_1136_0 | v_11693_0;
  assign v_1136_0 = v_1137_0 | v_11692_0;
  assign v_1137_0 = v_589_0 ? v_1138_0 : 3'h0;
  assign v_1139_0 = v_1140_0 | v_1141_0;
  assign v_1140_0 = v_589_0 | v_601_0;
  assign v_1141_0 = v_607_0 | v_26_0;
  assign v_1142_0 = v_1143_0 | v_11689_0;
  assign v_1143_0 = v_1144_0 | v_11688_0;
  assign v_1144_0 = v_589_0 ? v_1145_0 : 3'h0;
  assign v_1146_0 = v_1147_0 | v_1148_0;
  assign v_1147_0 = v_589_0 | v_601_0;
  assign v_1148_0 = v_607_0 | v_26_0;
  assign v_1149_0 = v_1150_0 | v_11685_0;
  assign v_1150_0 = v_1151_0 | v_11684_0;
  assign v_1151_0 = v_589_0 ? v_1152_0 : 3'h0;
  assign v_1153_0 = v_1154_0 | v_1155_0;
  assign v_1154_0 = v_589_0 | v_601_0;
  assign v_1155_0 = v_607_0 | v_26_0;
  assign v_1156_0 = v_1157_0 | v_11681_0;
  assign v_1157_0 = v_1158_0 | v_11680_0;
  assign v_1158_0 = v_589_0 ? v_1159_0 : 3'h0;
  assign v_1160_0 = v_1161_0 | v_1162_0;
  assign v_1161_0 = v_589_0 | v_601_0;
  assign v_1162_0 = v_607_0 | v_26_0;
  assign v_1163_0 = v_1164_0 | v_11677_0;
  assign v_1164_0 = v_1165_0 | v_11676_0;
  assign v_1165_0 = v_589_0 ? v_1166_0 : 3'h0;
  assign v_1167_0 = v_1168_0 | v_1169_0;
  assign v_1168_0 = v_589_0 | v_601_0;
  assign v_1169_0 = v_607_0 | v_26_0;
  assign v_1170_0 = v_1171_0 | v_11673_0;
  assign v_1171_0 = v_1172_0 | v_11672_0;
  assign v_1172_0 = v_589_0 ? v_1173_0 : 3'h0;
  assign v_1174_0 = v_1175_0 | v_1176_0;
  assign v_1175_0 = v_589_0 | v_601_0;
  assign v_1176_0 = v_607_0 | v_26_0;
  assign v_1177_0 = v_1178_0 | v_11669_0;
  assign v_1178_0 = v_1179_0 | v_11668_0;
  assign v_1179_0 = v_589_0 ? v_1180_0 : 3'h0;
  assign v_1181_0 = v_1182_0 | v_1183_0;
  assign v_1182_0 = v_589_0 | v_601_0;
  assign v_1183_0 = v_607_0 | v_26_0;
  assign v_1184_0 = v_1185_0 | v_11665_0;
  assign v_1185_0 = v_1186_0 | v_11664_0;
  assign v_1186_0 = v_589_0 ? v_1187_0 : 3'h0;
  assign v_1188_0 = v_1189_0 | v_1190_0;
  assign v_1189_0 = v_589_0 | v_601_0;
  assign v_1190_0 = v_607_0 | v_26_0;
  assign v_1191_0 = v_1192_0 | v_11661_0;
  assign v_1192_0 = v_1193_0 | v_11660_0;
  assign v_1193_0 = v_589_0 ? v_1194_0 : 3'h0;
  assign v_1195_0 = v_1196_0 | v_1197_0;
  assign v_1196_0 = v_589_0 | v_601_0;
  assign v_1197_0 = v_607_0 | v_26_0;
  assign v_1198_0 = v_1199_0 | v_11657_0;
  assign v_1199_0 = v_1200_0 | v_11656_0;
  assign v_1200_0 = v_589_0 ? v_1201_0 : 3'h0;
  assign v_1202_0 = v_1203_0 | v_1204_0;
  assign v_1203_0 = v_589_0 | v_601_0;
  assign v_1204_0 = v_607_0 | v_26_0;
  assign v_1205_0 = v_1206_0 | v_11653_0;
  assign v_1206_0 = v_1207_0 | v_11652_0;
  assign v_1207_0 = v_589_0 ? v_1208_0 : 3'h0;
  assign v_1209_0 = v_1210_0 | v_1211_0;
  assign v_1210_0 = v_589_0 | v_601_0;
  assign v_1211_0 = v_607_0 | v_26_0;
  assign v_1212_0 = v_1213_0 | v_11649_0;
  assign v_1213_0 = v_1214_0 | v_11648_0;
  assign v_1214_0 = v_589_0 ? v_1215_0 : 3'h0;
  assign v_1216_0 = v_1217_0 | v_1218_0;
  assign v_1217_0 = v_589_0 | v_601_0;
  assign v_1218_0 = v_607_0 | v_26_0;
  assign v_1219_0 = v_1220_0 | v_11645_0;
  assign v_1220_0 = v_1221_0 | v_11644_0;
  assign v_1221_0 = v_589_0 ? v_1222_0 : 3'h0;
  assign v_1223_0 = v_1224_0 | v_1225_0;
  assign v_1224_0 = v_589_0 | v_601_0;
  assign v_1225_0 = v_607_0 | v_26_0;
  assign v_1226_0 = v_1227_0 | v_11641_0;
  assign v_1227_0 = v_1228_0 | v_11640_0;
  assign v_1228_0 = v_589_0 ? v_1229_0 : 3'h0;
  assign v_1230_0 = v_1231_0 | v_1232_0;
  assign v_1231_0 = v_589_0 | v_601_0;
  assign v_1232_0 = v_607_0 | v_26_0;
  assign v_1233_0 = v_1234_0 | v_11637_0;
  assign v_1234_0 = v_1235_0 | v_11636_0;
  assign v_1235_0 = v_589_0 ? v_1236_0 : 3'h0;
  assign v_1237_0 = v_1238_0 | v_1239_0;
  assign v_1238_0 = v_589_0 | v_601_0;
  assign v_1239_0 = v_607_0 | v_26_0;
  assign v_1240_0 = v_1241_0 | v_11633_0;
  assign v_1241_0 = v_1242_0 | v_11632_0;
  assign v_1242_0 = v_589_0 ? v_1243_0 : 3'h0;
  assign v_1244_0 = v_1245_0 | v_1246_0;
  assign v_1245_0 = v_589_0 | v_601_0;
  assign v_1246_0 = v_607_0 | v_26_0;
  assign v_1247_0 = v_1248_0 | v_11629_0;
  assign v_1248_0 = v_1249_0 | v_11628_0;
  assign v_1249_0 = v_589_0 ? v_1250_0 : 3'h0;
  assign v_1251_0 = v_1252_0 | v_1253_0;
  assign v_1252_0 = v_589_0 | v_601_0;
  assign v_1253_0 = v_607_0 | v_26_0;
  assign v_1254_0 = v_1255_0 | v_11625_0;
  assign v_1255_0 = v_1256_0 | v_11624_0;
  assign v_1256_0 = v_589_0 ? v_1257_0 : 3'h0;
  assign v_1258_0 = v_1259_0 | v_1260_0;
  assign v_1259_0 = v_589_0 | v_601_0;
  assign v_1260_0 = v_607_0 | v_26_0;
  assign v_1261_0 = v_1262_0 | v_11621_0;
  assign v_1262_0 = v_1263_0 | v_11620_0;
  assign v_1263_0 = v_589_0 ? v_1264_0 : 3'h0;
  assign v_1265_0 = v_1266_0 | v_1267_0;
  assign v_1266_0 = v_589_0 | v_601_0;
  assign v_1267_0 = v_607_0 | v_26_0;
  assign v_1268_0 = v_1269_0 | v_11617_0;
  assign v_1269_0 = v_1270_0 | v_11616_0;
  assign v_1270_0 = v_589_0 ? v_1271_0 : 3'h0;
  assign v_1272_0 = v_1273_0 | v_1274_0;
  assign v_1273_0 = v_589_0 | v_601_0;
  assign v_1274_0 = v_607_0 | v_26_0;
  assign v_1275_0 = v_1276_0 | v_11613_0;
  assign v_1276_0 = v_1277_0 | v_11612_0;
  assign v_1277_0 = v_589_0 ? v_1278_0 : 3'h0;
  assign v_1279_0 = v_1280_0 | v_1281_0;
  assign v_1280_0 = v_589_0 | v_601_0;
  assign v_1281_0 = v_607_0 | v_26_0;
  assign v_1282_0 = v_1283_0 | v_11609_0;
  assign v_1283_0 = v_1284_0 | v_11608_0;
  assign v_1284_0 = v_589_0 ? v_1285_0 : 3'h0;
  assign v_1286_0 = v_1287_0 | v_1288_0;
  assign v_1287_0 = v_589_0 | v_601_0;
  assign v_1288_0 = v_607_0 | v_26_0;
  assign v_1289_0 = v_1290_0 | v_11605_0;
  assign v_1290_0 = v_1291_0 | v_11604_0;
  assign v_1291_0 = v_589_0 ? v_1292_0 : 3'h0;
  assign v_1293_0 = v_1294_0 | v_1295_0;
  assign v_1294_0 = v_589_0 | v_601_0;
  assign v_1295_0 = v_607_0 | v_26_0;
  assign v_1296_0 = v_1297_0 | v_11601_0;
  assign v_1297_0 = v_1298_0 | v_11600_0;
  assign v_1298_0 = v_589_0 ? v_1299_0 : 3'h0;
  assign v_1300_0 = v_1301_0 | v_1302_0;
  assign v_1301_0 = v_589_0 | v_601_0;
  assign v_1302_0 = v_607_0 | v_26_0;
  assign v_1303_0 = v_1304_0 | v_11597_0;
  assign v_1304_0 = v_1305_0 | v_11596_0;
  assign v_1305_0 = v_589_0 ? v_1306_0 : 3'h0;
  assign v_1307_0 = v_1308_0 | v_1309_0;
  assign v_1308_0 = v_589_0 | v_601_0;
  assign v_1309_0 = v_607_0 | v_26_0;
  assign v_1310_0 = v_1311_0 | v_11593_0;
  assign v_1311_0 = v_1312_0 | v_11592_0;
  assign v_1312_0 = v_589_0 ? v_1313_0 : 3'h0;
  assign v_1314_0 = v_1315_0 | v_1316_0;
  assign v_1315_0 = v_589_0 | v_601_0;
  assign v_1316_0 = v_607_0 | v_26_0;
  assign v_1317_0 = v_1318_0 | v_11589_0;
  assign v_1318_0 = v_1319_0 | v_11588_0;
  assign v_1319_0 = v_589_0 ? v_1320_0 : 3'h0;
  assign v_1321_0 = v_1322_0 | v_1323_0;
  assign v_1322_0 = v_589_0 | v_601_0;
  assign v_1323_0 = v_607_0 | v_26_0;
  assign v_1324_0 = v_1325_0 | v_11585_0;
  assign v_1325_0 = v_1326_0 | v_11584_0;
  assign v_1326_0 = v_589_0 ? v_1327_0 : 3'h0;
  assign v_1328_0 = v_1329_0 | v_1330_0;
  assign v_1329_0 = v_589_0 | v_601_0;
  assign v_1330_0 = v_607_0 | v_26_0;
  assign v_1331_0 = v_1332_0 | v_11581_0;
  assign v_1332_0 = v_1333_0 | v_11580_0;
  assign v_1333_0 = v_589_0 ? v_1334_0 : 3'h0;
  assign v_1335_0 = v_1336_0 | v_1337_0;
  assign v_1336_0 = v_589_0 | v_601_0;
  assign v_1337_0 = v_607_0 | v_26_0;
  assign v_1338_0 = v_1339_0 | v_11577_0;
  assign v_1339_0 = v_1340_0 | v_11576_0;
  assign v_1340_0 = v_589_0 ? v_1341_0 : 3'h0;
  assign v_1342_0 = v_1343_0 | v_1344_0;
  assign v_1343_0 = v_589_0 | v_601_0;
  assign v_1344_0 = v_607_0 | v_26_0;
  assign v_1345_0 = v_1346_0 | v_11573_0;
  assign v_1346_0 = v_1347_0 | v_11572_0;
  assign v_1347_0 = v_589_0 ? v_1348_0 : 3'h0;
  assign v_1349_0 = v_1350_0 | v_1351_0;
  assign v_1350_0 = v_589_0 | v_601_0;
  assign v_1351_0 = v_607_0 | v_26_0;
  assign v_1352_0 = v_1353_0 | v_11569_0;
  assign v_1353_0 = v_1354_0 | v_11568_0;
  assign v_1354_0 = v_589_0 ? v_1355_0 : 3'h0;
  assign v_1356_0 = v_1357_0 | v_1358_0;
  assign v_1357_0 = v_589_0 | v_601_0;
  assign v_1358_0 = v_607_0 | v_26_0;
  assign v_1359_0 = v_1360_0 | v_11565_0;
  assign v_1360_0 = v_1361_0 | v_11564_0;
  assign v_1361_0 = v_589_0 ? v_1362_0 : 3'h0;
  assign v_1363_0 = v_1364_0 | v_1365_0;
  assign v_1364_0 = v_589_0 | v_601_0;
  assign v_1365_0 = v_607_0 | v_26_0;
  assign v_1366_0 = v_1367_0 | v_11561_0;
  assign v_1367_0 = v_1368_0 | v_11560_0;
  assign v_1368_0 = v_589_0 ? v_1369_0 : 3'h0;
  assign v_1370_0 = v_1371_0 | v_1372_0;
  assign v_1371_0 = v_589_0 | v_601_0;
  assign v_1372_0 = v_607_0 | v_26_0;
  assign v_1373_0 = v_1374_0 | v_11557_0;
  assign v_1374_0 = v_1375_0 | v_11556_0;
  assign v_1375_0 = v_589_0 ? v_1376_0 : 3'h0;
  assign v_1377_0 = v_1378_0 | v_1379_0;
  assign v_1378_0 = v_589_0 | v_601_0;
  assign v_1379_0 = v_607_0 | v_26_0;
  assign v_1380_0 = v_1381_0 | v_11553_0;
  assign v_1381_0 = v_1382_0 | v_11552_0;
  assign v_1382_0 = v_589_0 ? v_1383_0 : 3'h0;
  assign v_1384_0 = v_1385_0 | v_1386_0;
  assign v_1385_0 = v_589_0 | v_601_0;
  assign v_1386_0 = v_607_0 | v_26_0;
  assign v_1387_0 = v_1388_0 | v_11549_0;
  assign v_1388_0 = v_1389_0 | v_11548_0;
  assign v_1389_0 = v_589_0 ? v_1390_0 : 3'h0;
  assign v_1391_0 = v_1392_0 | v_1393_0;
  assign v_1392_0 = v_589_0 | v_601_0;
  assign v_1393_0 = v_607_0 | v_26_0;
  assign v_1394_0 = v_1395_0 | v_11545_0;
  assign v_1395_0 = v_1396_0 | v_11544_0;
  assign v_1396_0 = v_589_0 ? v_1397_0 : 3'h0;
  assign v_1398_0 = v_1399_0 | v_1400_0;
  assign v_1399_0 = v_589_0 | v_601_0;
  assign v_1400_0 = v_607_0 | v_26_0;
  assign v_1401_0 = v_1402_0 | v_11541_0;
  assign v_1402_0 = v_1403_0 | v_11540_0;
  assign v_1403_0 = v_589_0 ? v_1404_0 : 3'h0;
  assign v_1405_0 = v_1406_0 | v_1407_0;
  assign v_1406_0 = v_589_0 | v_601_0;
  assign v_1407_0 = v_607_0 | v_26_0;
  assign v_1408_0 = v_1409_0 | v_11537_0;
  assign v_1409_0 = v_1410_0 | v_11536_0;
  assign v_1410_0 = v_589_0 ? v_1411_0 : 3'h0;
  assign v_1412_0 = v_1413_0 | v_1414_0;
  assign v_1413_0 = v_589_0 | v_601_0;
  assign v_1414_0 = v_607_0 | v_26_0;
  assign v_1415_0 = v_1416_0 | v_11533_0;
  assign v_1416_0 = v_1417_0 | v_11532_0;
  assign v_1417_0 = v_589_0 ? v_1418_0 : 3'h0;
  assign v_1419_0 = v_1420_0 | v_1421_0;
  assign v_1420_0 = v_589_0 | v_601_0;
  assign v_1421_0 = v_607_0 | v_26_0;
  assign v_1422_0 = v_1423_0 | v_11529_0;
  assign v_1423_0 = v_1424_0 | v_11528_0;
  assign v_1424_0 = v_589_0 ? v_1425_0 : 3'h0;
  assign v_1426_0 = v_1427_0 | v_1428_0;
  assign v_1427_0 = v_589_0 | v_601_0;
  assign v_1428_0 = v_607_0 | v_26_0;
  assign v_1429_0 = v_1430_0 | v_11525_0;
  assign v_1430_0 = v_1431_0 | v_11524_0;
  assign v_1431_0 = v_589_0 ? v_1432_0 : 3'h0;
  assign v_1433_0 = v_1434_0 | v_1435_0;
  assign v_1434_0 = v_589_0 | v_601_0;
  assign v_1435_0 = v_607_0 | v_26_0;
  assign v_1436_0 = v_1437_0 | v_11521_0;
  assign v_1437_0 = v_1438_0 | v_11520_0;
  assign v_1438_0 = v_589_0 ? v_1439_0 : 3'h0;
  assign v_1440_0 = v_1441_0 | v_1442_0;
  assign v_1441_0 = v_589_0 | v_601_0;
  assign v_1442_0 = v_607_0 | v_26_0;
  assign v_1443_0 = v_1444_0 | v_11517_0;
  assign v_1444_0 = v_1445_0 | v_11516_0;
  assign v_1445_0 = v_589_0 ? v_1446_0 : 3'h0;
  assign v_1447_0 = v_1448_0 | v_1449_0;
  assign v_1448_0 = v_589_0 | v_601_0;
  assign v_1449_0 = v_607_0 | v_26_0;
  assign v_1450_0 = v_1451_0 | v_11513_0;
  assign v_1451_0 = v_1452_0 | v_11512_0;
  assign v_1452_0 = v_589_0 ? v_1453_0 : 3'h0;
  assign v_1454_0 = v_1455_0 | v_1456_0;
  assign v_1455_0 = v_589_0 | v_601_0;
  assign v_1456_0 = v_607_0 | v_26_0;
  assign v_1457_0 = v_1458_0 | v_11509_0;
  assign v_1458_0 = v_1459_0 | v_11508_0;
  assign v_1459_0 = v_589_0 ? v_1460_0 : 3'h0;
  assign v_1461_0 = v_1462_0 | v_1463_0;
  assign v_1462_0 = v_589_0 | v_601_0;
  assign v_1463_0 = v_607_0 | v_26_0;
  assign v_1464_0 = v_1465_0 | v_11505_0;
  assign v_1465_0 = v_1466_0 | v_11504_0;
  assign v_1466_0 = v_589_0 ? v_1467_0 : 3'h0;
  assign v_1468_0 = v_1469_0 | v_1470_0;
  assign v_1469_0 = v_589_0 | v_601_0;
  assign v_1470_0 = v_607_0 | v_26_0;
  assign v_1471_0 = v_1472_0 | v_11501_0;
  assign v_1472_0 = v_1473_0 | v_11500_0;
  assign v_1473_0 = v_589_0 ? v_1474_0 : 3'h0;
  assign v_1475_0 = v_1476_0 | v_1477_0;
  assign v_1476_0 = v_589_0 | v_601_0;
  assign v_1477_0 = v_607_0 | v_26_0;
  assign v_1478_0 = v_1479_0 | v_11497_0;
  assign v_1479_0 = v_1480_0 | v_11496_0;
  assign v_1480_0 = v_589_0 ? v_1481_0 : 3'h0;
  assign v_1482_0 = v_1483_0 | v_1484_0;
  assign v_1483_0 = v_589_0 | v_601_0;
  assign v_1484_0 = v_607_0 | v_26_0;
  assign v_1485_0 = v_1486_0 | v_11493_0;
  assign v_1486_0 = v_1487_0 | v_11492_0;
  assign v_1487_0 = v_589_0 ? v_1488_0 : 3'h0;
  assign v_1489_0 = v_1490_0 | v_1491_0;
  assign v_1490_0 = v_589_0 | v_601_0;
  assign v_1491_0 = v_607_0 | v_26_0;
  assign v_1492_0 = v_1493_0 | v_11489_0;
  assign v_1493_0 = v_1494_0 | v_11488_0;
  assign v_1494_0 = v_589_0 ? v_1495_0 : 3'h0;
  assign v_1496_0 = v_1497_0 | v_1498_0;
  assign v_1497_0 = v_589_0 | v_601_0;
  assign v_1498_0 = v_607_0 | v_26_0;
  assign v_1499_0 = v_1500_0 | v_11485_0;
  assign v_1500_0 = v_1501_0 | v_11484_0;
  assign v_1501_0 = v_589_0 ? v_1502_0 : 3'h0;
  assign v_1503_0 = v_1504_0 | v_1505_0;
  assign v_1504_0 = v_589_0 | v_601_0;
  assign v_1505_0 = v_607_0 | v_26_0;
  assign v_1506_0 = v_1507_0 | v_11481_0;
  assign v_1507_0 = v_1508_0 | v_11480_0;
  assign v_1508_0 = v_589_0 ? v_1509_0 : 3'h0;
  assign v_1510_0 = v_1511_0 | v_1512_0;
  assign v_1511_0 = v_589_0 | v_601_0;
  assign v_1512_0 = v_607_0 | v_26_0;
  assign v_1513_0 = v_1514_0 | v_11477_0;
  assign v_1514_0 = v_1515_0 | v_11476_0;
  assign v_1515_0 = v_589_0 ? v_1516_0 : 3'h0;
  assign v_1517_0 = v_1518_0 | v_1519_0;
  assign v_1518_0 = v_589_0 | v_601_0;
  assign v_1519_0 = v_607_0 | v_26_0;
  assign v_1520_0 = v_1521_0 | v_11473_0;
  assign v_1521_0 = v_1522_0 | v_11472_0;
  assign v_1522_0 = v_589_0 ? v_1523_0 : 3'h0;
  assign v_1524_0 = v_1525_0 | v_1526_0;
  assign v_1525_0 = v_589_0 | v_601_0;
  assign v_1526_0 = v_607_0 | v_26_0;
  assign v_1527_0 = v_1528_0 | v_11469_0;
  assign v_1528_0 = v_1529_0 | v_11468_0;
  assign v_1529_0 = v_589_0 ? v_1530_0 : 3'h0;
  assign v_1531_0 = v_1532_0 | v_1533_0;
  assign v_1532_0 = v_589_0 | v_601_0;
  assign v_1533_0 = v_607_0 | v_26_0;
  assign v_1534_0 = v_1535_0 | v_11465_0;
  assign v_1535_0 = v_1536_0 | v_11464_0;
  assign v_1536_0 = v_589_0 ? v_1537_0 : 3'h0;
  assign v_1538_0 = v_1539_0 | v_1540_0;
  assign v_1539_0 = v_589_0 | v_601_0;
  assign v_1540_0 = v_607_0 | v_26_0;
  assign v_1541_0 = v_1542_0 | v_11461_0;
  assign v_1542_0 = v_1543_0 | v_11460_0;
  assign v_1543_0 = v_589_0 ? v_1544_0 : 3'h0;
  assign v_1545_0 = v_1546_0 | v_1547_0;
  assign v_1546_0 = v_589_0 | v_601_0;
  assign v_1547_0 = v_607_0 | v_26_0;
  assign v_1548_0 = v_1549_0 | v_11457_0;
  assign v_1549_0 = v_1550_0 | v_11456_0;
  assign v_1550_0 = v_589_0 ? v_1551_0 : 3'h0;
  assign v_1552_0 = v_1553_0 | v_1554_0;
  assign v_1553_0 = v_589_0 | v_601_0;
  assign v_1554_0 = v_607_0 | v_26_0;
  assign v_1555_0 = v_1556_0 | v_11453_0;
  assign v_1556_0 = v_1557_0 | v_11452_0;
  assign v_1557_0 = v_589_0 ? v_1558_0 : 3'h0;
  assign v_1559_0 = v_1560_0 | v_1561_0;
  assign v_1560_0 = v_589_0 | v_601_0;
  assign v_1561_0 = v_607_0 | v_26_0;
  assign v_1562_0 = v_1563_0 | v_11449_0;
  assign v_1563_0 = v_1564_0 | v_11448_0;
  assign v_1564_0 = v_589_0 ? v_1565_0 : 3'h0;
  assign v_1566_0 = v_1567_0 | v_1568_0;
  assign v_1567_0 = v_589_0 | v_601_0;
  assign v_1568_0 = v_607_0 | v_26_0;
  assign v_1569_0 = v_1570_0 | v_11445_0;
  assign v_1570_0 = v_1571_0 | v_11444_0;
  assign v_1571_0 = v_589_0 ? v_1572_0 : 3'h0;
  assign v_1573_0 = v_1574_0 | v_1575_0;
  assign v_1574_0 = v_589_0 | v_601_0;
  assign v_1575_0 = v_607_0 | v_26_0;
  assign v_1576_0 = v_1577_0 | v_11441_0;
  assign v_1577_0 = v_1578_0 | v_11440_0;
  assign v_1578_0 = v_589_0 ? v_1579_0 : 3'h0;
  assign v_1580_0 = v_1581_0 | v_1582_0;
  assign v_1581_0 = v_589_0 | v_601_0;
  assign v_1582_0 = v_607_0 | v_26_0;
  assign v_1583_0 = v_1584_0 | v_11437_0;
  assign v_1584_0 = v_1585_0 | v_11436_0;
  assign v_1585_0 = v_589_0 ? v_1586_0 : 3'h0;
  assign v_1587_0 = v_1588_0 | v_1589_0;
  assign v_1588_0 = v_589_0 | v_601_0;
  assign v_1589_0 = v_607_0 | v_26_0;
  assign v_1590_0 = v_1591_0 | v_11433_0;
  assign v_1591_0 = v_1592_0 | v_11432_0;
  assign v_1592_0 = v_589_0 ? v_1593_0 : 3'h0;
  assign v_1594_0 = v_1595_0 | v_1596_0;
  assign v_1595_0 = v_589_0 | v_601_0;
  assign v_1596_0 = v_607_0 | v_26_0;
  assign v_1597_0 = v_1598_0 | v_11429_0;
  assign v_1598_0 = v_1599_0 | v_11428_0;
  assign v_1599_0 = v_589_0 ? v_1600_0 : 3'h0;
  assign v_1601_0 = v_1602_0 | v_1603_0;
  assign v_1602_0 = v_589_0 | v_601_0;
  assign v_1603_0 = v_607_0 | v_26_0;
  assign v_1604_0 = v_1605_0 | v_11425_0;
  assign v_1605_0 = v_1606_0 | v_11424_0;
  assign v_1606_0 = v_589_0 ? v_1607_0 : 3'h0;
  assign v_1608_0 = v_1609_0 | v_1610_0;
  assign v_1609_0 = v_589_0 | v_601_0;
  assign v_1610_0 = v_607_0 | v_26_0;
  assign v_1611_0 = v_1612_0 | v_11421_0;
  assign v_1612_0 = v_1613_0 | v_11420_0;
  assign v_1613_0 = v_589_0 ? v_1614_0 : 3'h0;
  assign v_1615_0 = v_1616_0 | v_1617_0;
  assign v_1616_0 = v_589_0 | v_601_0;
  assign v_1617_0 = v_607_0 | v_26_0;
  assign v_1618_0 = v_1619_0 | v_11417_0;
  assign v_1619_0 = v_1620_0 | v_11416_0;
  assign v_1620_0 = v_589_0 ? v_1621_0 : 3'h0;
  assign v_1622_0 = v_1623_0 | v_1624_0;
  assign v_1623_0 = v_589_0 | v_601_0;
  assign v_1624_0 = v_607_0 | v_26_0;
  assign v_1625_0 = v_1626_0 | v_11413_0;
  assign v_1626_0 = v_1627_0 | v_11412_0;
  assign v_1627_0 = v_589_0 ? v_1628_0 : 3'h0;
  assign v_1629_0 = v_1630_0 | v_1631_0;
  assign v_1630_0 = v_589_0 | v_601_0;
  assign v_1631_0 = v_607_0 | v_26_0;
  assign v_1632_0 = v_1633_0 | v_11409_0;
  assign v_1633_0 = v_1634_0 | v_11408_0;
  assign v_1634_0 = v_589_0 ? v_1635_0 : 3'h0;
  assign v_1636_0 = v_1637_0 | v_1638_0;
  assign v_1637_0 = v_589_0 | v_601_0;
  assign v_1638_0 = v_607_0 | v_26_0;
  assign v_1639_0 = v_1640_0 | v_11405_0;
  assign v_1640_0 = v_1641_0 | v_11404_0;
  assign v_1641_0 = v_589_0 ? v_1642_0 : 3'h0;
  assign v_1643_0 = v_1644_0 | v_1645_0;
  assign v_1644_0 = v_589_0 | v_601_0;
  assign v_1645_0 = v_607_0 | v_26_0;
  assign v_1646_0 = v_1647_0 | v_11401_0;
  assign v_1647_0 = v_1648_0 | v_11400_0;
  assign v_1648_0 = v_589_0 ? v_1649_0 : 3'h0;
  assign v_1650_0 = v_1651_0 | v_1652_0;
  assign v_1651_0 = v_589_0 | v_601_0;
  assign v_1652_0 = v_607_0 | v_26_0;
  assign v_1653_0 = v_1654_0 | v_11397_0;
  assign v_1654_0 = v_1655_0 | v_11396_0;
  assign v_1655_0 = v_589_0 ? v_1656_0 : 3'h0;
  assign v_1657_0 = v_1658_0 | v_1659_0;
  assign v_1658_0 = v_589_0 | v_601_0;
  assign v_1659_0 = v_607_0 | v_26_0;
  assign v_1660_0 = v_1661_0 | v_11393_0;
  assign v_1661_0 = v_1662_0 | v_11392_0;
  assign v_1662_0 = v_589_0 ? v_1663_0 : 3'h0;
  assign v_1664_0 = v_1665_0 | v_1666_0;
  assign v_1665_0 = v_589_0 | v_601_0;
  assign v_1666_0 = v_607_0 | v_26_0;
  assign v_1667_0 = v_1668_0 | v_11389_0;
  assign v_1668_0 = v_1669_0 | v_11388_0;
  assign v_1669_0 = v_589_0 ? v_1670_0 : 3'h0;
  assign v_1671_0 = v_1672_0 | v_1673_0;
  assign v_1672_0 = v_589_0 | v_601_0;
  assign v_1673_0 = v_607_0 | v_26_0;
  assign v_1674_0 = v_1675_0 | v_11385_0;
  assign v_1675_0 = v_1676_0 | v_11384_0;
  assign v_1676_0 = v_589_0 ? v_1677_0 : 3'h0;
  assign v_1678_0 = v_1679_0 | v_1680_0;
  assign v_1679_0 = v_589_0 | v_601_0;
  assign v_1680_0 = v_607_0 | v_26_0;
  assign v_1681_0 = v_1682_0 | v_11381_0;
  assign v_1682_0 = v_1683_0 | v_11380_0;
  assign v_1683_0 = v_589_0 ? v_1684_0 : 3'h0;
  assign v_1685_0 = v_1686_0 | v_1687_0;
  assign v_1686_0 = v_589_0 | v_601_0;
  assign v_1687_0 = v_607_0 | v_26_0;
  assign v_1688_0 = v_1689_0 | v_11377_0;
  assign v_1689_0 = v_1690_0 | v_11376_0;
  assign v_1690_0 = v_589_0 ? v_1691_0 : 3'h0;
  assign v_1692_0 = v_1693_0 | v_1694_0;
  assign v_1693_0 = v_589_0 | v_601_0;
  assign v_1694_0 = v_607_0 | v_26_0;
  assign v_1695_0 = v_1696_0 | v_11373_0;
  assign v_1696_0 = v_1697_0 | v_11372_0;
  assign v_1697_0 = v_589_0 ? v_1698_0 : 3'h0;
  assign v_1699_0 = v_1700_0 | v_1701_0;
  assign v_1700_0 = v_589_0 | v_601_0;
  assign v_1701_0 = v_607_0 | v_26_0;
  assign v_1702_0 = v_1703_0 | v_11369_0;
  assign v_1703_0 = v_1704_0 | v_11368_0;
  assign v_1704_0 = v_589_0 ? v_1705_0 : 3'h0;
  assign v_1706_0 = v_1707_0 | v_1708_0;
  assign v_1707_0 = v_589_0 | v_601_0;
  assign v_1708_0 = v_607_0 | v_26_0;
  assign v_1709_0 = v_1710_0 | v_11365_0;
  assign v_1710_0 = v_1711_0 | v_11364_0;
  assign v_1711_0 = v_589_0 ? v_1712_0 : 3'h0;
  assign v_1713_0 = v_1714_0 | v_1715_0;
  assign v_1714_0 = v_589_0 | v_601_0;
  assign v_1715_0 = v_607_0 | v_26_0;
  assign v_1716_0 = v_1717_0 | v_11361_0;
  assign v_1717_0 = v_1718_0 | v_11360_0;
  assign v_1718_0 = v_589_0 ? v_1719_0 : 3'h0;
  assign v_1720_0 = v_1721_0 | v_1722_0;
  assign v_1721_0 = v_589_0 | v_601_0;
  assign v_1722_0 = v_607_0 | v_26_0;
  assign v_1723_0 = v_1724_0 | v_11357_0;
  assign v_1724_0 = v_1725_0 | v_11356_0;
  assign v_1725_0 = v_589_0 ? v_1726_0 : 3'h0;
  assign v_1727_0 = v_1728_0 | v_1729_0;
  assign v_1728_0 = v_589_0 | v_601_0;
  assign v_1729_0 = v_607_0 | v_26_0;
  assign v_1730_0 = v_1731_0 | v_11353_0;
  assign v_1731_0 = v_1732_0 | v_11352_0;
  assign v_1732_0 = v_589_0 ? v_1733_0 : 3'h0;
  assign v_1734_0 = v_1735_0 | v_1736_0;
  assign v_1735_0 = v_589_0 | v_601_0;
  assign v_1736_0 = v_607_0 | v_26_0;
  assign v_1737_0 = v_1738_0 | v_11349_0;
  assign v_1738_0 = v_1739_0 | v_11348_0;
  assign v_1739_0 = v_589_0 ? v_1740_0 : 3'h0;
  assign v_1741_0 = v_1742_0 | v_1743_0;
  assign v_1742_0 = v_589_0 | v_601_0;
  assign v_1743_0 = v_607_0 | v_26_0;
  assign v_1744_0 = v_1745_0 | v_11345_0;
  assign v_1745_0 = v_1746_0 | v_11344_0;
  assign v_1746_0 = v_589_0 ? v_1747_0 : 3'h0;
  assign v_1748_0 = v_1749_0 | v_1750_0;
  assign v_1749_0 = v_589_0 | v_601_0;
  assign v_1750_0 = v_607_0 | v_26_0;
  assign v_1751_0 = v_1752_0 | v_11341_0;
  assign v_1752_0 = v_1753_0 | v_11340_0;
  assign v_1753_0 = v_589_0 ? v_1754_0 : 3'h0;
  assign v_1755_0 = v_1756_0 | v_1757_0;
  assign v_1756_0 = v_589_0 | v_601_0;
  assign v_1757_0 = v_607_0 | v_26_0;
  assign v_1758_0 = v_1759_0 | v_11337_0;
  assign v_1759_0 = v_1760_0 | v_11336_0;
  assign v_1760_0 = v_589_0 ? v_1761_0 : 3'h0;
  assign v_1762_0 = v_1763_0 | v_1764_0;
  assign v_1763_0 = v_589_0 | v_601_0;
  assign v_1764_0 = v_607_0 | v_26_0;
  assign v_1765_0 = v_1766_0 | v_11333_0;
  assign v_1766_0 = v_1767_0 | v_11332_0;
  assign v_1767_0 = v_589_0 ? v_1768_0 : 3'h0;
  assign v_1769_0 = v_1770_0 | v_1771_0;
  assign v_1770_0 = v_589_0 | v_601_0;
  assign v_1771_0 = v_607_0 | v_26_0;
  assign v_1772_0 = v_1773_0 | v_11329_0;
  assign v_1773_0 = v_1774_0 | v_11328_0;
  assign v_1774_0 = v_589_0 ? v_1775_0 : 3'h0;
  assign v_1776_0 = v_1777_0 | v_1778_0;
  assign v_1777_0 = v_589_0 | v_601_0;
  assign v_1778_0 = v_607_0 | v_26_0;
  assign v_1779_0 = v_1780_0 | v_11325_0;
  assign v_1780_0 = v_1781_0 | v_11324_0;
  assign v_1781_0 = v_589_0 ? v_1782_0 : 3'h0;
  assign v_1783_0 = v_1784_0 | v_1785_0;
  assign v_1784_0 = v_589_0 | v_601_0;
  assign v_1785_0 = v_607_0 | v_26_0;
  assign v_1786_0 = v_1787_0 | v_11321_0;
  assign v_1787_0 = v_1788_0 | v_11320_0;
  assign v_1788_0 = v_589_0 ? v_1789_0 : 3'h0;
  assign v_1790_0 = v_1791_0 | v_1792_0;
  assign v_1791_0 = v_589_0 | v_601_0;
  assign v_1792_0 = v_607_0 | v_26_0;
  assign v_1793_0 = v_1794_0 | v_11317_0;
  assign v_1794_0 = v_1795_0 | v_11316_0;
  assign v_1795_0 = v_589_0 ? v_1796_0 : 3'h0;
  assign v_1797_0 = v_1798_0 | v_1799_0;
  assign v_1798_0 = v_589_0 | v_601_0;
  assign v_1799_0 = v_607_0 | v_26_0;
  assign v_1800_0 = v_1801_0 | v_11313_0;
  assign v_1801_0 = v_1802_0 | v_11312_0;
  assign v_1802_0 = v_589_0 ? v_1803_0 : 3'h0;
  assign v_1804_0 = v_1805_0 | v_1806_0;
  assign v_1805_0 = v_589_0 | v_601_0;
  assign v_1806_0 = v_607_0 | v_26_0;
  assign v_1807_0 = v_1808_0 | v_11309_0;
  assign v_1808_0 = v_1809_0 | v_11308_0;
  assign v_1809_0 = v_589_0 ? v_1810_0 : 3'h0;
  assign v_1811_0 = v_1812_0 | v_1813_0;
  assign v_1812_0 = v_589_0 | v_601_0;
  assign v_1813_0 = v_607_0 | v_26_0;
  assign v_1814_0 = v_1815_0 | v_11305_0;
  assign v_1815_0 = v_1816_0 | v_11304_0;
  assign v_1816_0 = v_589_0 ? v_1817_0 : 3'h0;
  assign v_1818_0 = v_1819_0 | v_1820_0;
  assign v_1819_0 = v_589_0 | v_601_0;
  assign v_1820_0 = v_607_0 | v_26_0;
  assign v_1821_0 = v_1822_0 | v_11301_0;
  assign v_1822_0 = v_1823_0 | v_11300_0;
  assign v_1823_0 = v_589_0 ? v_1824_0 : 3'h0;
  assign v_1825_0 = v_1826_0 | v_1827_0;
  assign v_1826_0 = v_589_0 | v_601_0;
  assign v_1827_0 = v_607_0 | v_26_0;
  assign v_1828_0 = v_1829_0 | v_11297_0;
  assign v_1829_0 = v_1830_0 | v_11296_0;
  assign v_1830_0 = v_589_0 ? v_1831_0 : 3'h0;
  assign v_1832_0 = v_1833_0 | v_1834_0;
  assign v_1833_0 = v_589_0 | v_601_0;
  assign v_1834_0 = v_607_0 | v_26_0;
  assign v_1835_0 = v_1836_0 | v_11293_0;
  assign v_1836_0 = v_1837_0 | v_11292_0;
  assign v_1837_0 = v_589_0 ? v_1838_0 : 3'h0;
  assign v_1839_0 = v_1840_0 | v_1841_0;
  assign v_1840_0 = v_589_0 | v_601_0;
  assign v_1841_0 = v_607_0 | v_26_0;
  assign v_1842_0 = v_1843_0 | v_11289_0;
  assign v_1843_0 = v_1844_0 | v_11288_0;
  assign v_1844_0 = v_589_0 ? v_1845_0 : 3'h0;
  assign v_1846_0 = v_1847_0 | v_1848_0;
  assign v_1847_0 = v_589_0 | v_601_0;
  assign v_1848_0 = v_607_0 | v_26_0;
  assign v_1849_0 = v_1850_0 | v_11285_0;
  assign v_1850_0 = v_1851_0 | v_11284_0;
  assign v_1851_0 = v_589_0 ? v_1852_0 : 3'h0;
  assign v_1853_0 = v_1854_0 | v_1855_0;
  assign v_1854_0 = v_589_0 | v_601_0;
  assign v_1855_0 = v_607_0 | v_26_0;
  assign v_1856_0 = v_1857_0 | v_11281_0;
  assign v_1857_0 = v_1858_0 | v_11280_0;
  assign v_1858_0 = v_589_0 ? v_1859_0 : 3'h0;
  assign v_1860_0 = v_1861_0 | v_1862_0;
  assign v_1861_0 = v_589_0 | v_601_0;
  assign v_1862_0 = v_607_0 | v_26_0;
  assign v_1863_0 = v_1864_0 | v_11277_0;
  assign v_1864_0 = v_1865_0 | v_11276_0;
  assign v_1865_0 = v_589_0 ? v_1866_0 : 3'h0;
  assign v_1867_0 = v_1868_0 | v_1869_0;
  assign v_1868_0 = v_589_0 | v_601_0;
  assign v_1869_0 = v_607_0 | v_26_0;
  assign v_1870_0 = v_1871_0 | v_11273_0;
  assign v_1871_0 = v_1872_0 | v_11272_0;
  assign v_1872_0 = v_589_0 ? v_1873_0 : 3'h0;
  assign v_1874_0 = v_1875_0 | v_1876_0;
  assign v_1875_0 = v_589_0 | v_601_0;
  assign v_1876_0 = v_607_0 | v_26_0;
  assign v_1877_0 = v_1878_0 | v_11269_0;
  assign v_1878_0 = v_1879_0 | v_11268_0;
  assign v_1879_0 = v_589_0 ? v_1880_0 : 3'h0;
  assign v_1881_0 = v_1882_0 | v_1883_0;
  assign v_1882_0 = v_589_0 | v_601_0;
  assign v_1883_0 = v_607_0 | v_26_0;
  assign v_1884_0 = v_1885_0 | v_11265_0;
  assign v_1885_0 = v_1886_0 | v_11264_0;
  assign v_1886_0 = v_589_0 ? v_1887_0 : 3'h0;
  assign v_1888_0 = v_1889_0 | v_1890_0;
  assign v_1889_0 = v_589_0 | v_601_0;
  assign v_1890_0 = v_607_0 | v_26_0;
  assign v_1891_0 = v_1892_0 | v_11261_0;
  assign v_1892_0 = v_1893_0 | v_11260_0;
  assign v_1893_0 = v_589_0 ? v_1894_0 : 3'h0;
  assign v_1895_0 = v_1896_0 | v_1897_0;
  assign v_1896_0 = v_589_0 | v_601_0;
  assign v_1897_0 = v_607_0 | v_26_0;
  assign v_1898_0 = v_1899_0 | v_11257_0;
  assign v_1899_0 = v_1900_0 | v_11256_0;
  assign v_1900_0 = v_589_0 ? v_1901_0 : 3'h0;
  assign v_1902_0 = v_1903_0 | v_1904_0;
  assign v_1903_0 = v_589_0 | v_601_0;
  assign v_1904_0 = v_607_0 | v_26_0;
  assign v_1905_0 = v_1906_0 | v_11253_0;
  assign v_1906_0 = v_1907_0 | v_11252_0;
  assign v_1907_0 = v_589_0 ? v_1908_0 : 3'h0;
  assign v_1909_0 = v_1910_0 | v_1911_0;
  assign v_1910_0 = v_589_0 | v_601_0;
  assign v_1911_0 = v_607_0 | v_26_0;
  assign v_1912_0 = v_1913_0 | v_11249_0;
  assign v_1913_0 = v_1914_0 | v_11248_0;
  assign v_1914_0 = v_589_0 ? v_1915_0 : 3'h0;
  assign v_1916_0 = v_1917_0 | v_1918_0;
  assign v_1917_0 = v_589_0 | v_601_0;
  assign v_1918_0 = v_607_0 | v_26_0;
  assign v_1919_0 = v_1920_0 | v_11245_0;
  assign v_1920_0 = v_1921_0 | v_11244_0;
  assign v_1921_0 = v_589_0 ? v_1922_0 : 3'h0;
  assign v_1923_0 = v_1924_0 | v_1925_0;
  assign v_1924_0 = v_589_0 | v_601_0;
  assign v_1925_0 = v_607_0 | v_26_0;
  assign v_1926_0 = v_1927_0 | v_11241_0;
  assign v_1927_0 = v_1928_0 | v_11240_0;
  assign v_1928_0 = v_589_0 ? v_1929_0 : 3'h0;
  assign v_1930_0 = v_1931_0 | v_1932_0;
  assign v_1931_0 = v_589_0 | v_601_0;
  assign v_1932_0 = v_607_0 | v_26_0;
  assign v_1933_0 = v_1934_0 | v_11237_0;
  assign v_1934_0 = v_1935_0 | v_11236_0;
  assign v_1935_0 = v_589_0 ? v_1936_0 : 3'h0;
  assign v_1937_0 = v_1938_0 | v_1939_0;
  assign v_1938_0 = v_589_0 | v_601_0;
  assign v_1939_0 = v_607_0 | v_26_0;
  assign v_1940_0 = v_1941_0 | v_11233_0;
  assign v_1941_0 = v_1942_0 | v_11232_0;
  assign v_1942_0 = v_589_0 ? v_1943_0 : 3'h0;
  assign v_1944_0 = v_1945_0 | v_1946_0;
  assign v_1945_0 = v_589_0 | v_601_0;
  assign v_1946_0 = v_607_0 | v_26_0;
  assign v_1947_0 = v_1948_0 | v_11229_0;
  assign v_1948_0 = v_1949_0 | v_11228_0;
  assign v_1949_0 = v_589_0 ? v_1950_0 : 3'h0;
  assign v_1951_0 = v_1952_0 | v_1953_0;
  assign v_1952_0 = v_589_0 | v_601_0;
  assign v_1953_0 = v_607_0 | v_26_0;
  assign v_1954_0 = v_1955_0 | v_11225_0;
  assign v_1955_0 = v_1956_0 | v_11224_0;
  assign v_1956_0 = v_589_0 ? v_1957_0 : 3'h0;
  assign v_1958_0 = v_1959_0 | v_1960_0;
  assign v_1959_0 = v_589_0 | v_601_0;
  assign v_1960_0 = v_607_0 | v_26_0;
  assign v_1961_0 = v_1962_0 | v_11221_0;
  assign v_1962_0 = v_1963_0 | v_11220_0;
  assign v_1963_0 = v_589_0 ? v_1964_0 : 3'h0;
  assign v_1965_0 = v_1966_0 | v_1967_0;
  assign v_1966_0 = v_589_0 | v_601_0;
  assign v_1967_0 = v_607_0 | v_26_0;
  assign v_1968_0 = v_1969_0 | v_11217_0;
  assign v_1969_0 = v_1970_0 | v_11216_0;
  assign v_1970_0 = v_589_0 ? v_1971_0 : 3'h0;
  assign v_1972_0 = v_1973_0 | v_1974_0;
  assign v_1973_0 = v_589_0 | v_601_0;
  assign v_1974_0 = v_607_0 | v_26_0;
  assign v_1975_0 = v_1976_0 | v_11213_0;
  assign v_1976_0 = v_1977_0 | v_11212_0;
  assign v_1977_0 = v_589_0 ? v_1978_0 : 3'h0;
  assign v_1979_0 = v_1980_0 | v_1981_0;
  assign v_1980_0 = v_589_0 | v_601_0;
  assign v_1981_0 = v_607_0 | v_26_0;
  assign v_1982_0 = v_1983_0 | v_11209_0;
  assign v_1983_0 = v_1984_0 | v_11208_0;
  assign v_1984_0 = v_589_0 ? v_1985_0 : 3'h0;
  assign v_1986_0 = v_1987_0 | v_1988_0;
  assign v_1987_0 = v_589_0 | v_601_0;
  assign v_1988_0 = v_607_0 | v_26_0;
  assign v_1989_0 = v_1990_0 | v_11205_0;
  assign v_1990_0 = v_1991_0 | v_11204_0;
  assign v_1991_0 = v_589_0 ? v_1992_0 : 3'h0;
  assign v_1993_0 = v_1994_0 | v_1995_0;
  assign v_1994_0 = v_589_0 | v_601_0;
  assign v_1995_0 = v_607_0 | v_26_0;
  assign v_1996_0 = v_1997_0 | v_11201_0;
  assign v_1997_0 = v_1998_0 | v_11200_0;
  assign v_1998_0 = v_589_0 ? v_1999_0 : 3'h0;
  assign v_2000_0 = v_2001_0 | v_2002_0;
  assign v_2001_0 = v_589_0 | v_601_0;
  assign v_2002_0 = v_607_0 | v_26_0;
  assign v_2003_0 = v_2004_0 | v_11197_0;
  assign v_2004_0 = v_2005_0 | v_11196_0;
  assign v_2005_0 = v_589_0 ? v_2006_0 : 3'h0;
  assign v_2007_0 = v_2008_0 | v_2009_0;
  assign v_2008_0 = v_589_0 | v_601_0;
  assign v_2009_0 = v_607_0 | v_26_0;
  assign v_2010_0 = v_2011_0 | v_11193_0;
  assign v_2011_0 = v_2012_0 | v_11192_0;
  assign v_2012_0 = v_589_0 ? v_2013_0 : 3'h0;
  assign v_2014_0 = v_2015_0 | v_2016_0;
  assign v_2015_0 = v_589_0 | v_601_0;
  assign v_2016_0 = v_607_0 | v_26_0;
  assign v_2017_0 = v_2018_0 | v_11189_0;
  assign v_2018_0 = v_2019_0 | v_11188_0;
  assign v_2019_0 = v_589_0 ? v_2020_0 : 3'h0;
  assign v_2021_0 = v_2022_0 | v_2023_0;
  assign v_2022_0 = v_589_0 | v_601_0;
  assign v_2023_0 = v_607_0 | v_26_0;
  assign v_2024_0 = v_2025_0 | v_11185_0;
  assign v_2025_0 = v_2026_0 | v_11184_0;
  assign v_2026_0 = v_589_0 ? v_2027_0 : 3'h0;
  assign v_2028_0 = v_2029_0 | v_2030_0;
  assign v_2029_0 = v_589_0 | v_601_0;
  assign v_2030_0 = v_607_0 | v_26_0;
  assign v_2031_0 = v_2032_0 | v_11181_0;
  assign v_2032_0 = v_2033_0 | v_11180_0;
  assign v_2033_0 = v_589_0 ? v_2034_0 : 3'h0;
  assign v_2035_0 = v_2036_0 | v_2037_0;
  assign v_2036_0 = v_589_0 | v_601_0;
  assign v_2037_0 = v_607_0 | v_26_0;
  assign v_2038_0 = v_2039_0 | v_11177_0;
  assign v_2039_0 = v_2040_0 | v_11176_0;
  assign v_2040_0 = v_589_0 ? v_2041_0 : 3'h0;
  assign v_2042_0 = v_2043_0 | v_2044_0;
  assign v_2043_0 = v_589_0 | v_601_0;
  assign v_2044_0 = v_607_0 | v_26_0;
  assign v_2045_0 = v_2046_0 | v_11173_0;
  assign v_2046_0 = v_2047_0 | v_11172_0;
  assign v_2047_0 = v_589_0 ? v_2048_0 : 3'h0;
  assign v_2049_0 = v_2050_0 | v_2051_0;
  assign v_2050_0 = v_589_0 | v_601_0;
  assign v_2051_0 = v_607_0 | v_26_0;
  assign v_2052_0 = v_2053_0 | v_11169_0;
  assign v_2053_0 = v_2054_0 | v_11168_0;
  assign v_2054_0 = v_589_0 ? v_2055_0 : 3'h0;
  assign v_2056_0 = v_2057_0 | v_2058_0;
  assign v_2057_0 = v_589_0 | v_601_0;
  assign v_2058_0 = v_607_0 | v_26_0;
  assign v_2059_0 = v_2060_0 | v_11165_0;
  assign v_2060_0 = v_2061_0 | v_11164_0;
  assign v_2061_0 = v_589_0 ? v_2062_0 : 3'h0;
  assign v_2063_0 = v_2064_0 | v_2065_0;
  assign v_2064_0 = v_589_0 | v_601_0;
  assign v_2065_0 = v_607_0 | v_26_0;
  assign v_2066_0 = v_2067_0 | v_11161_0;
  assign v_2067_0 = v_2068_0 | v_11160_0;
  assign v_2068_0 = v_589_0 ? v_2069_0 : 3'h0;
  assign v_2070_0 = v_2071_0 | v_2072_0;
  assign v_2071_0 = v_589_0 | v_601_0;
  assign v_2072_0 = v_607_0 | v_26_0;
  assign v_2073_0 = v_2074_0 | v_11157_0;
  assign v_2074_0 = v_2075_0 | v_11156_0;
  assign v_2075_0 = v_589_0 ? v_2076_0 : 3'h0;
  assign v_2077_0 = v_2078_0 | v_2079_0;
  assign v_2078_0 = v_589_0 | v_601_0;
  assign v_2079_0 = v_607_0 | v_26_0;
  assign v_2080_0 = v_2081_0 | v_11153_0;
  assign v_2081_0 = v_2082_0 | v_11152_0;
  assign v_2082_0 = v_589_0 ? v_2083_0 : 3'h0;
  assign v_2084_0 = v_2085_0 | v_2086_0;
  assign v_2085_0 = v_589_0 | v_601_0;
  assign v_2086_0 = v_607_0 | v_26_0;
  assign v_2087_0 = v_2088_0 | v_11149_0;
  assign v_2088_0 = v_2089_0 | v_11148_0;
  assign v_2089_0 = v_589_0 ? v_2090_0 : 3'h0;
  assign v_2091_0 = v_2092_0 | v_2093_0;
  assign v_2092_0 = v_589_0 | v_601_0;
  assign v_2093_0 = v_607_0 | v_26_0;
  assign v_2094_0 = v_2095_0 | v_11145_0;
  assign v_2095_0 = v_2096_0 | v_11144_0;
  assign v_2096_0 = v_589_0 ? v_2097_0 : 3'h0;
  assign v_2098_0 = v_2099_0 | v_2100_0;
  assign v_2099_0 = v_589_0 | v_601_0;
  assign v_2100_0 = v_607_0 | v_26_0;
  assign v_2101_0 = v_2102_0 | v_11141_0;
  assign v_2102_0 = v_2103_0 | v_11140_0;
  assign v_2103_0 = v_589_0 ? v_2104_0 : 3'h0;
  assign v_2105_0 = v_2106_0 | v_2107_0;
  assign v_2106_0 = v_589_0 | v_601_0;
  assign v_2107_0 = v_607_0 | v_26_0;
  assign v_2108_0 = v_2109_0 | v_11137_0;
  assign v_2109_0 = v_2110_0 | v_11136_0;
  assign v_2110_0 = v_589_0 ? v_2111_0 : 3'h0;
  assign v_2112_0 = v_2113_0 | v_2114_0;
  assign v_2113_0 = v_589_0 | v_601_0;
  assign v_2114_0 = v_607_0 | v_26_0;
  assign v_2115_0 = v_2116_0 | v_11133_0;
  assign v_2116_0 = v_2117_0 | v_11132_0;
  assign v_2117_0 = v_589_0 ? v_2118_0 : 3'h0;
  assign v_2119_0 = v_2120_0 | v_2121_0;
  assign v_2120_0 = v_589_0 | v_601_0;
  assign v_2121_0 = v_607_0 | v_26_0;
  assign v_2122_0 = v_2123_0 | v_11129_0;
  assign v_2123_0 = v_2124_0 | v_11128_0;
  assign v_2124_0 = v_589_0 ? v_2125_0 : 3'h0;
  assign v_2126_0 = v_2127_0 | v_2128_0;
  assign v_2127_0 = v_589_0 | v_601_0;
  assign v_2128_0 = v_607_0 | v_26_0;
  assign v_2129_0 = v_2130_0 | v_11125_0;
  assign v_2130_0 = v_2131_0 | v_11124_0;
  assign v_2131_0 = v_589_0 ? v_2132_0 : 3'h0;
  assign v_2133_0 = v_2134_0 | v_2135_0;
  assign v_2134_0 = v_589_0 | v_601_0;
  assign v_2135_0 = v_607_0 | v_26_0;
  assign v_2136_0 = v_2137_0 | v_11121_0;
  assign v_2137_0 = v_2138_0 | v_11120_0;
  assign v_2138_0 = v_589_0 ? v_2139_0 : 3'h0;
  assign v_2140_0 = v_2141_0 | v_2142_0;
  assign v_2141_0 = v_589_0 | v_601_0;
  assign v_2142_0 = v_607_0 | v_26_0;
  assign v_2143_0 = v_2144_0 | v_11117_0;
  assign v_2144_0 = v_2145_0 | v_11116_0;
  assign v_2145_0 = v_589_0 ? v_2146_0 : 3'h0;
  assign v_2147_0 = v_2148_0 | v_2149_0;
  assign v_2148_0 = v_589_0 | v_601_0;
  assign v_2149_0 = v_607_0 | v_26_0;
  assign v_2150_0 = v_2151_0 | v_11113_0;
  assign v_2151_0 = v_2152_0 | v_11112_0;
  assign v_2152_0 = v_589_0 ? v_2153_0 : 3'h0;
  assign v_2154_0 = v_2155_0 | v_2156_0;
  assign v_2155_0 = v_589_0 | v_601_0;
  assign v_2156_0 = v_607_0 | v_26_0;
  assign v_2157_0 = v_2158_0 | v_11109_0;
  assign v_2158_0 = v_2159_0 | v_11108_0;
  assign v_2159_0 = v_589_0 ? v_2160_0 : 3'h0;
  assign v_2161_0 = v_2162_0 | v_2163_0;
  assign v_2162_0 = v_589_0 | v_601_0;
  assign v_2163_0 = v_607_0 | v_26_0;
  assign v_2164_0 = v_2165_0 | v_11105_0;
  assign v_2165_0 = v_2166_0 | v_11104_0;
  assign v_2166_0 = v_589_0 ? v_2167_0 : 3'h0;
  assign v_2168_0 = v_2169_0 | v_2170_0;
  assign v_2169_0 = v_589_0 | v_601_0;
  assign v_2170_0 = v_607_0 | v_26_0;
  assign v_2171_0 = v_2172_0 | v_11101_0;
  assign v_2172_0 = v_2173_0 | v_11100_0;
  assign v_2173_0 = v_589_0 ? v_2174_0 : 3'h0;
  assign v_2175_0 = v_2176_0 | v_2177_0;
  assign v_2176_0 = v_589_0 | v_601_0;
  assign v_2177_0 = v_607_0 | v_26_0;
  assign v_2178_0 = v_2179_0 | v_11097_0;
  assign v_2179_0 = v_2180_0 | v_11096_0;
  assign v_2180_0 = v_589_0 ? v_2181_0 : 3'h0;
  assign v_2182_0 = v_2183_0 | v_2184_0;
  assign v_2183_0 = v_589_0 | v_601_0;
  assign v_2184_0 = v_607_0 | v_26_0;
  assign v_2185_0 = v_2186_0 | v_11093_0;
  assign v_2186_0 = v_2187_0 | v_11092_0;
  assign v_2187_0 = v_589_0 ? v_2188_0 : 3'h0;
  assign v_2189_0 = v_2190_0 | v_2191_0;
  assign v_2190_0 = v_589_0 | v_601_0;
  assign v_2191_0 = v_607_0 | v_26_0;
  assign v_2192_0 = v_2193_0 | v_11089_0;
  assign v_2193_0 = v_2194_0 | v_11088_0;
  assign v_2194_0 = v_589_0 ? v_2195_0 : 3'h0;
  assign v_2196_0 = v_2197_0 | v_2198_0;
  assign v_2197_0 = v_589_0 | v_601_0;
  assign v_2198_0 = v_607_0 | v_26_0;
  assign v_2199_0 = v_2200_0 | v_11085_0;
  assign v_2200_0 = v_2201_0 | v_11084_0;
  assign v_2201_0 = v_589_0 ? v_2202_0 : 3'h0;
  assign v_2203_0 = v_2204_0 | v_2205_0;
  assign v_2204_0 = v_589_0 | v_601_0;
  assign v_2205_0 = v_607_0 | v_26_0;
  assign v_2206_0 = v_2207_0 | v_11081_0;
  assign v_2207_0 = v_2208_0 | v_11080_0;
  assign v_2208_0 = v_589_0 ? v_2209_0 : 3'h0;
  assign v_2210_0 = v_2211_0 | v_2212_0;
  assign v_2211_0 = v_589_0 | v_601_0;
  assign v_2212_0 = v_607_0 | v_26_0;
  assign v_2213_0 = v_2214_0 | v_11077_0;
  assign v_2214_0 = v_2215_0 | v_11076_0;
  assign v_2215_0 = v_589_0 ? v_2216_0 : 3'h0;
  assign v_2217_0 = v_2218_0 | v_2219_0;
  assign v_2218_0 = v_589_0 | v_601_0;
  assign v_2219_0 = v_607_0 | v_26_0;
  assign v_2220_0 = v_2221_0 | v_11073_0;
  assign v_2221_0 = v_2222_0 | v_11072_0;
  assign v_2222_0 = v_589_0 ? v_2223_0 : 3'h0;
  assign v_2224_0 = v_2225_0 | v_2226_0;
  assign v_2225_0 = v_589_0 | v_601_0;
  assign v_2226_0 = v_607_0 | v_26_0;
  assign v_2227_0 = v_2228_0 | v_11069_0;
  assign v_2228_0 = v_2229_0 | v_11068_0;
  assign v_2229_0 = v_589_0 ? v_2230_0 : 3'h0;
  assign v_2231_0 = v_2232_0 | v_2233_0;
  assign v_2232_0 = v_589_0 | v_601_0;
  assign v_2233_0 = v_607_0 | v_26_0;
  assign v_2234_0 = v_2235_0 | v_11065_0;
  assign v_2235_0 = v_2236_0 | v_11064_0;
  assign v_2236_0 = v_589_0 ? v_2237_0 : 3'h0;
  assign v_2238_0 = v_2239_0 | v_2240_0;
  assign v_2239_0 = v_589_0 | v_601_0;
  assign v_2240_0 = v_607_0 | v_26_0;
  assign v_2241_0 = v_2242_0 | v_11061_0;
  assign v_2242_0 = v_2243_0 | v_11060_0;
  assign v_2243_0 = v_589_0 ? v_2244_0 : 3'h0;
  assign v_2245_0 = v_2246_0 | v_2247_0;
  assign v_2246_0 = v_589_0 | v_601_0;
  assign v_2247_0 = v_607_0 | v_26_0;
  assign v_2248_0 = v_2249_0 | v_11057_0;
  assign v_2249_0 = v_2250_0 | v_11056_0;
  assign v_2250_0 = v_589_0 ? v_2251_0 : 3'h0;
  assign v_2252_0 = v_2253_0 | v_2254_0;
  assign v_2253_0 = v_589_0 | v_601_0;
  assign v_2254_0 = v_607_0 | v_26_0;
  assign v_2255_0 = v_2256_0 | v_11053_0;
  assign v_2256_0 = v_2257_0 | v_11052_0;
  assign v_2257_0 = v_589_0 ? v_2258_0 : 3'h0;
  assign v_2259_0 = v_2260_0 | v_2261_0;
  assign v_2260_0 = v_589_0 | v_601_0;
  assign v_2261_0 = v_607_0 | v_26_0;
  assign v_2262_0 = v_2263_0 | v_11049_0;
  assign v_2263_0 = v_2264_0 | v_11048_0;
  assign v_2264_0 = v_589_0 ? v_2265_0 : 3'h0;
  assign v_2266_0 = v_2267_0 | v_2268_0;
  assign v_2267_0 = v_589_0 | v_601_0;
  assign v_2268_0 = v_607_0 | v_26_0;
  assign v_2269_0 = v_2270_0 | v_11045_0;
  assign v_2270_0 = v_2271_0 | v_11044_0;
  assign v_2271_0 = v_589_0 ? v_2272_0 : 3'h0;
  assign v_2273_0 = v_2274_0 | v_2275_0;
  assign v_2274_0 = v_589_0 | v_601_0;
  assign v_2275_0 = v_607_0 | v_26_0;
  assign v_2276_0 = v_2277_0 | v_11041_0;
  assign v_2277_0 = v_2278_0 | v_11040_0;
  assign v_2278_0 = v_589_0 ? v_2279_0 : 3'h0;
  assign v_2280_0 = v_2281_0 | v_2282_0;
  assign v_2281_0 = v_589_0 | v_601_0;
  assign v_2282_0 = v_607_0 | v_26_0;
  assign v_2283_0 = v_2284_0 | v_11037_0;
  assign v_2284_0 = v_2285_0 | v_11036_0;
  assign v_2285_0 = v_589_0 ? v_2286_0 : 3'h0;
  assign v_2287_0 = v_2288_0 | v_2289_0;
  assign v_2288_0 = v_589_0 | v_601_0;
  assign v_2289_0 = v_607_0 | v_26_0;
  assign v_2290_0 = v_2291_0 | v_11033_0;
  assign v_2291_0 = v_2292_0 | v_11032_0;
  assign v_2292_0 = v_589_0 ? v_2293_0 : 3'h0;
  assign v_2294_0 = v_2295_0 | v_2296_0;
  assign v_2295_0 = v_589_0 | v_601_0;
  assign v_2296_0 = v_607_0 | v_26_0;
  assign v_2297_0 = v_2298_0 | v_11029_0;
  assign v_2298_0 = v_2299_0 | v_11028_0;
  assign v_2299_0 = v_589_0 ? v_2300_0 : 3'h0;
  assign v_2301_0 = v_2302_0 | v_2303_0;
  assign v_2302_0 = v_589_0 | v_601_0;
  assign v_2303_0 = v_607_0 | v_26_0;
  assign v_2304_0 = v_2305_0 | v_11025_0;
  assign v_2305_0 = v_2306_0 | v_11024_0;
  assign v_2306_0 = v_589_0 ? v_2307_0 : 3'h0;
  assign v_2308_0 = v_2309_0 | v_2310_0;
  assign v_2309_0 = v_589_0 | v_601_0;
  assign v_2310_0 = v_607_0 | v_26_0;
  assign v_2311_0 = v_2312_0 | v_11021_0;
  assign v_2312_0 = v_2313_0 | v_11020_0;
  assign v_2313_0 = v_589_0 ? v_2314_0 : 3'h0;
  assign v_2315_0 = v_2316_0 | v_2317_0;
  assign v_2316_0 = v_589_0 | v_601_0;
  assign v_2317_0 = v_607_0 | v_26_0;
  assign v_2318_0 = v_2319_0 | v_11017_0;
  assign v_2319_0 = v_2320_0 | v_11016_0;
  assign v_2320_0 = v_589_0 ? v_2321_0 : 3'h0;
  assign v_2322_0 = v_2323_0 | v_2324_0;
  assign v_2323_0 = v_589_0 | v_601_0;
  assign v_2324_0 = v_607_0 | v_26_0;
  assign v_2325_0 = v_2326_0 | v_11013_0;
  assign v_2326_0 = v_2327_0 | v_11012_0;
  assign v_2327_0 = v_589_0 ? v_2328_0 : 3'h0;
  assign v_2329_0 = v_2330_0 | v_2331_0;
  assign v_2330_0 = v_589_0 | v_601_0;
  assign v_2331_0 = v_607_0 | v_26_0;
  assign v_2332_0 = v_2333_0 | v_11009_0;
  assign v_2333_0 = v_2334_0 | v_11008_0;
  assign v_2334_0 = v_589_0 ? v_2335_0 : 3'h0;
  assign v_2336_0 = v_2337_0 | v_2338_0;
  assign v_2337_0 = v_589_0 | v_601_0;
  assign v_2338_0 = v_607_0 | v_26_0;
  assign v_2339_0 = v_2340_0 | v_11005_0;
  assign v_2340_0 = v_2341_0 | v_11004_0;
  assign v_2341_0 = v_589_0 ? v_2342_0 : 3'h0;
  assign v_2343_0 = v_2344_0 | v_2345_0;
  assign v_2344_0 = v_589_0 | v_601_0;
  assign v_2345_0 = v_607_0 | v_26_0;
  assign v_2346_0 = v_2347_0 | v_11001_0;
  assign v_2347_0 = v_2348_0 | v_11000_0;
  assign v_2348_0 = v_589_0 ? v_2349_0 : 3'h0;
  assign v_2350_0 = v_2351_0 | v_2352_0;
  assign v_2351_0 = v_589_0 | v_601_0;
  assign v_2352_0 = v_607_0 | v_26_0;
  assign v_2353_0 = v_2354_0 | v_10997_0;
  assign v_2354_0 = v_2355_0 | v_10996_0;
  assign v_2355_0 = v_589_0 ? v_2356_0 : 3'h0;
  assign v_2357_0 = v_2358_0 | v_2359_0;
  assign v_2358_0 = v_589_0 | v_601_0;
  assign v_2359_0 = v_607_0 | v_26_0;
  assign v_2360_0 = v_2361_0 | v_10993_0;
  assign v_2361_0 = v_2362_0 | v_10992_0;
  assign v_2362_0 = v_589_0 ? v_2363_0 : 3'h0;
  assign v_2364_0 = v_2365_0 | v_2366_0;
  assign v_2365_0 = v_589_0 | v_601_0;
  assign v_2366_0 = v_607_0 | v_26_0;
  assign v_2367_0 = v_2368_0 | v_10989_0;
  assign v_2368_0 = v_2369_0 | v_10988_0;
  assign v_2369_0 = v_589_0 ? v_2370_0 : 3'h0;
  assign v_2371_0 = v_2372_0 | v_2373_0;
  assign v_2372_0 = v_589_0 | v_601_0;
  assign v_2373_0 = v_607_0 | v_26_0;
  assign v_2374_0 = v_2375_0 | v_10985_0;
  assign v_2375_0 = v_2376_0 | v_10984_0;
  assign v_2376_0 = v_589_0 ? v_2377_0 : 3'h0;
  assign v_2378_0 = v_2379_0 | v_2380_0;
  assign v_2379_0 = v_589_0 | v_601_0;
  assign v_2380_0 = v_607_0 | v_26_0;
  assign v_2381_0 = v_2382_0 | v_10981_0;
  assign v_2382_0 = v_2383_0 | v_10980_0;
  assign v_2383_0 = v_589_0 ? v_2384_0 : 3'h0;
  assign v_2385_0 = v_2386_0 | v_2387_0;
  assign v_2386_0 = v_589_0 | v_601_0;
  assign v_2387_0 = v_607_0 | v_26_0;
  assign v_2388_0 = v_2389_0 | v_10977_0;
  assign v_2389_0 = v_2390_0 | v_10976_0;
  assign v_2390_0 = v_589_0 ? v_2391_0 : 3'h0;
  assign v_2392_0 = v_2393_0 | v_2394_0;
  assign v_2393_0 = v_589_0 | v_601_0;
  assign v_2394_0 = v_607_0 | v_26_0;
  assign v_2395_0 = v_2396_0 | v_10973_0;
  assign v_2396_0 = v_2397_0 | v_10972_0;
  assign v_2397_0 = v_589_0 ? v_2398_0 : 3'h0;
  assign v_2399_0 = v_2400_0 | v_2401_0;
  assign v_2400_0 = v_589_0 | v_601_0;
  assign v_2401_0 = v_607_0 | v_26_0;
  assign v_2402_0 = v_2403_0 | v_10969_0;
  assign v_2403_0 = v_2404_0 | v_10968_0;
  assign v_2404_0 = v_589_0 ? v_2405_0 : 3'h0;
  assign v_2406_0 = v_2407_0 | v_2408_0;
  assign v_2407_0 = v_589_0 | v_601_0;
  assign v_2408_0 = v_607_0 | v_26_0;
  assign v_2409_0 = v_2410_0 | v_10965_0;
  assign v_2410_0 = v_2411_0 | v_10964_0;
  assign v_2411_0 = v_589_0 ? v_2412_0 : 3'h0;
  assign v_2413_0 = v_2414_0 | v_2415_0;
  assign v_2414_0 = v_589_0 | v_601_0;
  assign v_2415_0 = v_607_0 | v_26_0;
  assign v_2416_0 = v_2417_0 | v_10961_0;
  assign v_2417_0 = v_2418_0 | v_10960_0;
  assign v_2418_0 = v_589_0 ? v_2419_0 : 3'h0;
  assign v_2420_0 = v_2421_0 | v_2422_0;
  assign v_2421_0 = v_589_0 | v_601_0;
  assign v_2422_0 = v_607_0 | v_26_0;
  assign v_2423_0 = v_2424_0 | v_10957_0;
  assign v_2424_0 = v_2425_0 | v_10956_0;
  assign v_2425_0 = v_589_0 ? v_2426_0 : 3'h0;
  assign v_2427_0 = v_2428_0 | v_2429_0;
  assign v_2428_0 = v_589_0 | v_601_0;
  assign v_2429_0 = v_607_0 | v_26_0;
  assign v_2430_0 = v_2431_0 | v_10953_0;
  assign v_2431_0 = v_2432_0 | v_10952_0;
  assign v_2432_0 = v_589_0 ? v_2433_0 : 3'h0;
  assign v_2434_0 = v_2435_0 | v_2436_0;
  assign v_2435_0 = v_589_0 | v_601_0;
  assign v_2436_0 = v_607_0 | v_26_0;
  assign v_2437_0 = v_2438_0 | v_10949_0;
  assign v_2438_0 = v_2439_0 | v_10948_0;
  assign v_2439_0 = v_589_0 ? v_2440_0 : 3'h0;
  assign v_2441_0 = v_2442_0 | v_2443_0;
  assign v_2442_0 = v_589_0 | v_601_0;
  assign v_2443_0 = v_607_0 | v_26_0;
  assign v_2444_0 = v_2445_0 | v_10945_0;
  assign v_2445_0 = v_2446_0 | v_10944_0;
  assign v_2446_0 = v_589_0 ? v_2447_0 : 3'h0;
  assign v_2448_0 = v_2449_0 | v_2450_0;
  assign v_2449_0 = v_589_0 | v_601_0;
  assign v_2450_0 = v_607_0 | v_26_0;
  assign v_2451_0 = v_2452_0 | v_10941_0;
  assign v_2452_0 = v_2453_0 | v_10940_0;
  assign v_2453_0 = v_589_0 ? v_2454_0 : 3'h0;
  assign v_2455_0 = v_2456_0 | v_2457_0;
  assign v_2456_0 = v_589_0 | v_601_0;
  assign v_2457_0 = v_607_0 | v_26_0;
  assign v_2458_0 = v_2459_0 | v_10937_0;
  assign v_2459_0 = v_2460_0 | v_10936_0;
  assign v_2460_0 = v_589_0 ? v_2461_0 : 3'h0;
  assign v_2462_0 = v_2463_0 | v_2464_0;
  assign v_2463_0 = v_589_0 | v_601_0;
  assign v_2464_0 = v_607_0 | v_26_0;
  assign v_2465_0 = v_2466_0 | v_10933_0;
  assign v_2466_0 = v_2467_0 | v_10932_0;
  assign v_2467_0 = v_589_0 ? v_2468_0 : 3'h0;
  assign v_2469_0 = v_2470_0 | v_2471_0;
  assign v_2470_0 = v_589_0 | v_601_0;
  assign v_2471_0 = v_607_0 | v_26_0;
  assign v_2472_0 = v_2473_0 | v_10929_0;
  assign v_2473_0 = v_2474_0 | v_10928_0;
  assign v_2474_0 = v_589_0 ? v_2475_0 : 3'h0;
  assign v_2476_0 = v_2477_0 | v_2478_0;
  assign v_2477_0 = v_589_0 | v_601_0;
  assign v_2478_0 = v_607_0 | v_26_0;
  assign v_2479_0 = v_2480_0 | v_10925_0;
  assign v_2480_0 = v_2481_0 | v_10924_0;
  assign v_2481_0 = v_589_0 ? v_2482_0 : 3'h0;
  assign v_2483_0 = v_2484_0 | v_2485_0;
  assign v_2484_0 = v_589_0 | v_601_0;
  assign v_2485_0 = v_607_0 | v_26_0;
  assign v_2486_0 = v_2487_0 | v_10921_0;
  assign v_2487_0 = v_2488_0 | v_10920_0;
  assign v_2488_0 = v_589_0 ? v_2489_0 : 3'h0;
  assign v_2490_0 = v_2491_0 | v_2492_0;
  assign v_2491_0 = v_589_0 | v_601_0;
  assign v_2492_0 = v_607_0 | v_26_0;
  assign v_2493_0 = v_2494_0 | v_10917_0;
  assign v_2494_0 = v_2495_0 | v_10916_0;
  assign v_2495_0 = v_589_0 ? v_2496_0 : 3'h0;
  assign v_2497_0 = v_2498_0 | v_2499_0;
  assign v_2498_0 = v_589_0 | v_601_0;
  assign v_2499_0 = v_607_0 | v_26_0;
  assign v_2500_0 = v_2501_0 | v_10913_0;
  assign v_2501_0 = v_2502_0 | v_10912_0;
  assign v_2502_0 = v_589_0 ? v_2503_0 : 3'h0;
  assign v_2504_0 = v_2505_0 | v_2506_0;
  assign v_2505_0 = v_589_0 | v_601_0;
  assign v_2506_0 = v_607_0 | v_26_0;
  assign v_2507_0 = v_2508_0 | v_10909_0;
  assign v_2508_0 = v_2509_0 | v_10908_0;
  assign v_2509_0 = v_589_0 ? v_2510_0 : 3'h0;
  assign v_2511_0 = v_2512_0 | v_2513_0;
  assign v_2512_0 = v_589_0 | v_601_0;
  assign v_2513_0 = v_607_0 | v_26_0;
  assign v_2514_0 = v_2515_0 | v_10905_0;
  assign v_2515_0 = v_2516_0 | v_10904_0;
  assign v_2516_0 = v_589_0 ? v_2517_0 : 3'h0;
  assign v_2518_0 = v_2519_0 | v_2520_0;
  assign v_2519_0 = v_589_0 | v_601_0;
  assign v_2520_0 = v_607_0 | v_26_0;
  assign v_2521_0 = v_2522_0 | v_10901_0;
  assign v_2522_0 = v_2523_0 | v_10900_0;
  assign v_2523_0 = v_589_0 ? v_2524_0 : 3'h0;
  assign v_2525_0 = v_2526_0 | v_2527_0;
  assign v_2526_0 = v_589_0 | v_601_0;
  assign v_2527_0 = v_607_0 | v_26_0;
  assign v_2528_0 = v_2529_0 | v_10897_0;
  assign v_2529_0 = v_2530_0 | v_10896_0;
  assign v_2530_0 = v_589_0 ? v_2531_0 : 3'h0;
  assign v_2532_0 = v_2533_0 | v_2534_0;
  assign v_2533_0 = v_589_0 | v_601_0;
  assign v_2534_0 = v_607_0 | v_26_0;
  assign v_2535_0 = v_2536_0 | v_10893_0;
  assign v_2536_0 = v_2537_0 | v_10892_0;
  assign v_2537_0 = v_589_0 ? v_2538_0 : 3'h0;
  assign v_2539_0 = v_2540_0 | v_2541_0;
  assign v_2540_0 = v_589_0 | v_601_0;
  assign v_2541_0 = v_607_0 | v_26_0;
  assign v_2542_0 = v_2543_0 | v_10889_0;
  assign v_2543_0 = v_2544_0 | v_10888_0;
  assign v_2544_0 = v_589_0 ? v_2545_0 : 3'h0;
  assign v_2546_0 = v_2547_0 | v_2548_0;
  assign v_2547_0 = v_589_0 | v_601_0;
  assign v_2548_0 = v_607_0 | v_26_0;
  assign v_2549_0 = v_2550_0 | v_10885_0;
  assign v_2550_0 = v_2551_0 | v_10884_0;
  assign v_2551_0 = v_589_0 ? v_2552_0 : 3'h0;
  assign v_2553_0 = v_2554_0 | v_2555_0;
  assign v_2554_0 = v_589_0 | v_601_0;
  assign v_2555_0 = v_607_0 | v_26_0;
  assign v_2556_0 = v_2557_0 | v_10881_0;
  assign v_2557_0 = v_2558_0 | v_10880_0;
  assign v_2558_0 = v_589_0 ? v_2559_0 : 3'h0;
  assign v_2560_0 = v_2561_0 | v_2562_0;
  assign v_2561_0 = v_589_0 | v_601_0;
  assign v_2562_0 = v_607_0 | v_26_0;
  assign v_2563_0 = v_2564_0 | v_10877_0;
  assign v_2564_0 = v_2565_0 | v_10876_0;
  assign v_2565_0 = v_589_0 ? v_2566_0 : 3'h0;
  assign v_2567_0 = v_2568_0 | v_2569_0;
  assign v_2568_0 = v_589_0 | v_601_0;
  assign v_2569_0 = v_607_0 | v_26_0;
  assign v_2570_0 = v_2571_0 | v_10873_0;
  assign v_2571_0 = v_2572_0 | v_10872_0;
  assign v_2572_0 = v_589_0 ? v_2573_0 : 3'h0;
  assign v_2574_0 = v_2575_0 | v_2576_0;
  assign v_2575_0 = v_589_0 | v_601_0;
  assign v_2576_0 = v_607_0 | v_26_0;
  assign v_2577_0 = v_2578_0 | v_10869_0;
  assign v_2578_0 = v_2579_0 | v_10868_0;
  assign v_2579_0 = v_589_0 ? v_2580_0 : 3'h0;
  assign v_2581_0 = v_2582_0 | v_2583_0;
  assign v_2582_0 = v_589_0 | v_601_0;
  assign v_2583_0 = v_607_0 | v_26_0;
  assign v_2584_0 = v_2585_0 | v_10865_0;
  assign v_2585_0 = v_2586_0 | v_10864_0;
  assign v_2586_0 = v_589_0 ? v_2587_0 : 3'h0;
  assign v_2588_0 = v_2589_0 | v_2590_0;
  assign v_2589_0 = v_589_0 | v_601_0;
  assign v_2590_0 = v_607_0 | v_26_0;
  assign v_2591_0 = v_2592_0 | v_10861_0;
  assign v_2592_0 = v_2593_0 | v_10860_0;
  assign v_2593_0 = v_589_0 ? v_2594_0 : 3'h0;
  assign v_2595_0 = v_2596_0 | v_2597_0;
  assign v_2596_0 = v_589_0 | v_601_0;
  assign v_2597_0 = v_607_0 | v_26_0;
  assign v_2598_0 = v_2599_0 | v_10857_0;
  assign v_2599_0 = v_2600_0 | v_10856_0;
  assign v_2600_0 = v_589_0 ? v_2601_0 : 3'h0;
  assign v_2602_0 = v_2603_0 | v_2604_0;
  assign v_2603_0 = v_589_0 | v_601_0;
  assign v_2604_0 = v_607_0 | v_26_0;
  assign v_2605_0 = v_2606_0 | v_10853_0;
  assign v_2606_0 = v_2607_0 | v_10852_0;
  assign v_2607_0 = v_589_0 ? v_2608_0 : 3'h0;
  assign v_2609_0 = v_2610_0 | v_2611_0;
  assign v_2610_0 = v_589_0 | v_601_0;
  assign v_2611_0 = v_607_0 | v_26_0;
  assign v_2612_0 = v_2613_0 | v_10849_0;
  assign v_2613_0 = v_2614_0 | v_10848_0;
  assign v_2614_0 = v_589_0 ? v_2615_0 : 3'h0;
  assign v_2616_0 = v_2617_0 | v_2618_0;
  assign v_2617_0 = v_589_0 | v_601_0;
  assign v_2618_0 = v_607_0 | v_26_0;
  assign v_2619_0 = v_2620_0 | v_10845_0;
  assign v_2620_0 = v_2621_0 | v_10844_0;
  assign v_2621_0 = v_589_0 ? v_2622_0 : 3'h0;
  assign v_2623_0 = v_2624_0 | v_2625_0;
  assign v_2624_0 = v_589_0 | v_601_0;
  assign v_2625_0 = v_607_0 | v_26_0;
  assign v_2626_0 = v_2627_0 | v_10841_0;
  assign v_2627_0 = v_2628_0 | v_10840_0;
  assign v_2628_0 = v_589_0 ? v_2629_0 : 3'h0;
  assign v_2630_0 = v_2631_0 | v_2632_0;
  assign v_2631_0 = v_589_0 | v_601_0;
  assign v_2632_0 = v_607_0 | v_26_0;
  assign v_2633_0 = v_2634_0 | v_10837_0;
  assign v_2634_0 = v_2635_0 | v_10836_0;
  assign v_2635_0 = v_589_0 ? v_2636_0 : 3'h0;
  assign v_2637_0 = v_2638_0 | v_2639_0;
  assign v_2638_0 = v_589_0 | v_601_0;
  assign v_2639_0 = v_607_0 | v_26_0;
  assign v_2640_0 = v_2641_0 | v_10833_0;
  assign v_2641_0 = v_2642_0 | v_10832_0;
  assign v_2642_0 = v_589_0 ? v_2643_0 : 3'h0;
  assign v_2644_0 = v_2645_0 | v_2646_0;
  assign v_2645_0 = v_589_0 | v_601_0;
  assign v_2646_0 = v_607_0 | v_26_0;
  assign v_2647_0 = v_2648_0 | v_10829_0;
  assign v_2648_0 = v_2649_0 | v_10828_0;
  assign v_2649_0 = v_589_0 ? v_2650_0 : 3'h0;
  assign v_2651_0 = v_2652_0 | v_2653_0;
  assign v_2652_0 = v_589_0 | v_601_0;
  assign v_2653_0 = v_607_0 | v_26_0;
  assign v_2654_0 = v_2655_0 | v_10825_0;
  assign v_2655_0 = v_2656_0 | v_10824_0;
  assign v_2656_0 = v_589_0 ? v_2657_0 : 3'h0;
  assign v_2658_0 = v_2659_0 | v_2660_0;
  assign v_2659_0 = v_589_0 | v_601_0;
  assign v_2660_0 = v_607_0 | v_26_0;
  assign v_2661_0 = v_2662_0 | v_10821_0;
  assign v_2662_0 = v_2663_0 | v_10820_0;
  assign v_2663_0 = v_589_0 ? v_2664_0 : 3'h0;
  assign v_2665_0 = v_2666_0 | v_2667_0;
  assign v_2666_0 = v_589_0 | v_601_0;
  assign v_2667_0 = v_607_0 | v_26_0;
  assign v_2668_0 = v_2669_0 | v_10817_0;
  assign v_2669_0 = v_2670_0 | v_10816_0;
  assign v_2670_0 = v_589_0 ? v_2671_0 : 3'h0;
  assign v_2672_0 = v_2673_0 | v_2674_0;
  assign v_2673_0 = v_589_0 | v_601_0;
  assign v_2674_0 = v_607_0 | v_26_0;
  assign v_2675_0 = v_2676_0 | v_10813_0;
  assign v_2676_0 = v_2677_0 | v_10812_0;
  assign v_2677_0 = v_589_0 ? v_2678_0 : 3'h0;
  assign v_2679_0 = v_2680_0 | v_2681_0;
  assign v_2680_0 = v_589_0 | v_601_0;
  assign v_2681_0 = v_607_0 | v_26_0;
  assign v_2682_0 = v_2683_0 | v_10809_0;
  assign v_2683_0 = v_2684_0 | v_10808_0;
  assign v_2684_0 = v_589_0 ? v_2685_0 : 3'h0;
  assign v_2686_0 = v_2687_0 | v_2688_0;
  assign v_2687_0 = v_589_0 | v_601_0;
  assign v_2688_0 = v_607_0 | v_26_0;
  assign v_2689_0 = v_2690_0 | v_10805_0;
  assign v_2690_0 = v_2691_0 | v_10804_0;
  assign v_2691_0 = v_589_0 ? v_2692_0 : 3'h0;
  assign v_2693_0 = v_2694_0 | v_2695_0;
  assign v_2694_0 = v_589_0 | v_601_0;
  assign v_2695_0 = v_607_0 | v_26_0;
  assign v_2696_0 = v_2697_0 | v_10801_0;
  assign v_2697_0 = v_2698_0 | v_10800_0;
  assign v_2698_0 = v_589_0 ? v_2699_0 : 3'h0;
  assign v_2700_0 = v_2701_0 | v_2702_0;
  assign v_2701_0 = v_589_0 | v_601_0;
  assign v_2702_0 = v_607_0 | v_26_0;
  assign v_2703_0 = v_2704_0 | v_10797_0;
  assign v_2704_0 = v_2705_0 | v_10796_0;
  assign v_2705_0 = v_589_0 ? v_2706_0 : 3'h0;
  assign v_2707_0 = v_2708_0 | v_2709_0;
  assign v_2708_0 = v_589_0 | v_601_0;
  assign v_2709_0 = v_607_0 | v_26_0;
  assign v_2710_0 = v_2711_0 | v_10793_0;
  assign v_2711_0 = v_2712_0 | v_10792_0;
  assign v_2712_0 = v_589_0 ? v_2713_0 : 3'h0;
  assign v_2714_0 = v_2715_0 | v_2716_0;
  assign v_2715_0 = v_589_0 | v_601_0;
  assign v_2716_0 = v_607_0 | v_26_0;
  assign v_2717_0 = v_2718_0 | v_10789_0;
  assign v_2718_0 = v_2719_0 | v_10788_0;
  assign v_2719_0 = v_589_0 ? v_2720_0 : 3'h0;
  assign v_2721_0 = v_2722_0 | v_2723_0;
  assign v_2722_0 = v_589_0 | v_601_0;
  assign v_2723_0 = v_607_0 | v_26_0;
  assign v_2724_0 = v_2725_0 | v_10785_0;
  assign v_2725_0 = v_2726_0 | v_10784_0;
  assign v_2726_0 = v_589_0 ? v_2727_0 : 3'h0;
  assign v_2728_0 = v_2729_0 | v_2730_0;
  assign v_2729_0 = v_589_0 | v_601_0;
  assign v_2730_0 = v_607_0 | v_26_0;
  assign v_2731_0 = v_2732_0 | v_10781_0;
  assign v_2732_0 = v_2733_0 | v_10780_0;
  assign v_2733_0 = v_589_0 ? v_2734_0 : 3'h0;
  assign v_2735_0 = v_2736_0 | v_2737_0;
  assign v_2736_0 = v_589_0 | v_601_0;
  assign v_2737_0 = v_607_0 | v_26_0;
  assign v_2738_0 = v_2739_0 | v_10777_0;
  assign v_2739_0 = v_2740_0 | v_10776_0;
  assign v_2740_0 = v_589_0 ? v_2741_0 : 3'h0;
  assign v_2742_0 = v_2743_0 | v_2744_0;
  assign v_2743_0 = v_589_0 | v_601_0;
  assign v_2744_0 = v_607_0 | v_26_0;
  assign v_2745_0 = v_2746_0 | v_10773_0;
  assign v_2746_0 = v_2747_0 | v_10772_0;
  assign v_2747_0 = v_589_0 ? v_2748_0 : 3'h0;
  assign v_2749_0 = v_2750_0 | v_2751_0;
  assign v_2750_0 = v_589_0 | v_601_0;
  assign v_2751_0 = v_607_0 | v_26_0;
  assign v_2752_0 = v_2753_0 | v_10769_0;
  assign v_2753_0 = v_2754_0 | v_10768_0;
  assign v_2754_0 = v_589_0 ? v_2755_0 : 3'h0;
  assign v_2756_0 = v_2757_0 | v_2758_0;
  assign v_2757_0 = v_589_0 | v_601_0;
  assign v_2758_0 = v_607_0 | v_26_0;
  assign v_2759_0 = v_2760_0 | v_10765_0;
  assign v_2760_0 = v_2761_0 | v_10764_0;
  assign v_2761_0 = v_589_0 ? v_2762_0 : 3'h0;
  assign v_2763_0 = v_2764_0 | v_2765_0;
  assign v_2764_0 = v_589_0 | v_601_0;
  assign v_2765_0 = v_607_0 | v_26_0;
  assign v_2766_0 = v_2767_0 | v_10761_0;
  assign v_2767_0 = v_2768_0 | v_10760_0;
  assign v_2768_0 = v_589_0 ? v_2769_0 : 3'h0;
  assign v_2770_0 = v_2771_0 | v_2772_0;
  assign v_2771_0 = v_589_0 | v_601_0;
  assign v_2772_0 = v_607_0 | v_26_0;
  assign v_2773_0 = v_2774_0 | v_10757_0;
  assign v_2774_0 = v_2775_0 | v_10756_0;
  assign v_2775_0 = v_589_0 ? v_2776_0 : 3'h0;
  assign v_2777_0 = v_2778_0 | v_2779_0;
  assign v_2778_0 = v_589_0 | v_601_0;
  assign v_2779_0 = v_607_0 | v_26_0;
  assign v_2780_0 = v_2781_0 | v_10753_0;
  assign v_2781_0 = v_2782_0 | v_10752_0;
  assign v_2782_0 = v_589_0 ? v_2783_0 : 3'h0;
  assign v_2784_0 = v_2785_0 | v_2786_0;
  assign v_2785_0 = v_589_0 | v_601_0;
  assign v_2786_0 = v_607_0 | v_26_0;
  assign v_2787_0 = v_2788_0 | v_10749_0;
  assign v_2788_0 = v_2789_0 | v_10748_0;
  assign v_2789_0 = v_589_0 ? v_2790_0 : 3'h0;
  assign v_2791_0 = v_2792_0 | v_2793_0;
  assign v_2792_0 = v_589_0 | v_601_0;
  assign v_2793_0 = v_607_0 | v_26_0;
  assign v_2794_0 = v_2795_0 | v_10745_0;
  assign v_2795_0 = v_2796_0 | v_10744_0;
  assign v_2796_0 = v_589_0 ? v_2797_0 : 3'h0;
  assign v_2798_0 = v_2799_0 | v_2800_0;
  assign v_2799_0 = v_589_0 | v_601_0;
  assign v_2800_0 = v_607_0 | v_26_0;
  assign v_2801_0 = v_2802_0 | v_10741_0;
  assign v_2802_0 = v_2803_0 | v_10740_0;
  assign v_2803_0 = v_589_0 ? v_2804_0 : 3'h0;
  assign v_2805_0 = v_2806_0 | v_2807_0;
  assign v_2806_0 = v_589_0 | v_601_0;
  assign v_2807_0 = v_607_0 | v_26_0;
  assign v_2808_0 = v_2809_0 | v_10737_0;
  assign v_2809_0 = v_2810_0 | v_10736_0;
  assign v_2810_0 = v_589_0 ? v_2811_0 : 3'h0;
  assign v_2812_0 = v_2813_0 | v_2814_0;
  assign v_2813_0 = v_589_0 | v_601_0;
  assign v_2814_0 = v_607_0 | v_26_0;
  assign v_2815_0 = v_2816_0 | v_10733_0;
  assign v_2816_0 = v_2817_0 | v_10732_0;
  assign v_2817_0 = v_589_0 ? v_2818_0 : 3'h0;
  assign v_2819_0 = v_2820_0 | v_2821_0;
  assign v_2820_0 = v_589_0 | v_601_0;
  assign v_2821_0 = v_607_0 | v_26_0;
  assign v_2822_0 = v_2823_0 | v_10729_0;
  assign v_2823_0 = v_2824_0 | v_10728_0;
  assign v_2824_0 = v_589_0 ? v_2825_0 : 3'h0;
  assign v_2826_0 = v_2827_0 | v_2828_0;
  assign v_2827_0 = v_589_0 | v_601_0;
  assign v_2828_0 = v_607_0 | v_26_0;
  assign v_2829_0 = v_2830_0 | v_10725_0;
  assign v_2830_0 = v_2831_0 | v_10724_0;
  assign v_2831_0 = v_589_0 ? v_2832_0 : 3'h0;
  assign v_2833_0 = v_2834_0 | v_2835_0;
  assign v_2834_0 = v_589_0 | v_601_0;
  assign v_2835_0 = v_607_0 | v_26_0;
  assign v_2836_0 = v_2837_0 | v_10721_0;
  assign v_2837_0 = v_2838_0 | v_10720_0;
  assign v_2838_0 = v_589_0 ? v_2839_0 : 3'h0;
  assign v_2840_0 = v_2841_0 | v_2842_0;
  assign v_2841_0 = v_589_0 | v_601_0;
  assign v_2842_0 = v_607_0 | v_26_0;
  assign v_2843_0 = v_2844_0 | v_10717_0;
  assign v_2844_0 = v_2845_0 | v_10716_0;
  assign v_2845_0 = v_589_0 ? v_2846_0 : 3'h0;
  assign v_2847_0 = v_2848_0 | v_2849_0;
  assign v_2848_0 = v_589_0 | v_601_0;
  assign v_2849_0 = v_607_0 | v_26_0;
  assign v_2850_0 = v_2851_0 | v_10713_0;
  assign v_2851_0 = v_2852_0 | v_10712_0;
  assign v_2852_0 = v_589_0 ? v_2853_0 : 3'h0;
  assign v_2854_0 = v_2855_0 | v_2856_0;
  assign v_2855_0 = v_589_0 | v_601_0;
  assign v_2856_0 = v_607_0 | v_26_0;
  assign v_2857_0 = v_2858_0 | v_10709_0;
  assign v_2858_0 = v_2859_0 | v_10708_0;
  assign v_2859_0 = v_589_0 ? v_2860_0 : 3'h0;
  assign v_2861_0 = v_2862_0 | v_2863_0;
  assign v_2862_0 = v_589_0 | v_601_0;
  assign v_2863_0 = v_607_0 | v_26_0;
  assign v_2864_0 = v_2865_0 | v_10705_0;
  assign v_2865_0 = v_2866_0 | v_10704_0;
  assign v_2866_0 = v_589_0 ? v_2867_0 : 3'h0;
  assign v_2868_0 = v_2869_0 | v_2870_0;
  assign v_2869_0 = v_589_0 | v_601_0;
  assign v_2870_0 = v_607_0 | v_26_0;
  assign v_2871_0 = v_2872_0 | v_10701_0;
  assign v_2872_0 = v_2873_0 | v_10700_0;
  assign v_2873_0 = v_589_0 ? v_2874_0 : 3'h0;
  assign v_2875_0 = v_2876_0 | v_2877_0;
  assign v_2876_0 = v_589_0 | v_601_0;
  assign v_2877_0 = v_607_0 | v_26_0;
  assign v_2878_0 = v_2879_0 | v_10697_0;
  assign v_2879_0 = v_2880_0 | v_10696_0;
  assign v_2880_0 = v_589_0 ? v_2881_0 : 3'h0;
  assign v_2882_0 = v_2883_0 | v_2884_0;
  assign v_2883_0 = v_589_0 | v_601_0;
  assign v_2884_0 = v_607_0 | v_26_0;
  assign v_2885_0 = v_2886_0 | v_10693_0;
  assign v_2886_0 = v_2887_0 | v_10692_0;
  assign v_2887_0 = v_589_0 ? v_2888_0 : 3'h0;
  assign v_2889_0 = v_2890_0 | v_2891_0;
  assign v_2890_0 = v_589_0 | v_601_0;
  assign v_2891_0 = v_607_0 | v_26_0;
  assign v_2892_0 = v_2893_0 | v_10689_0;
  assign v_2893_0 = v_2894_0 | v_10688_0;
  assign v_2894_0 = v_589_0 ? v_2895_0 : 3'h0;
  assign v_2896_0 = v_2897_0 | v_2898_0;
  assign v_2897_0 = v_589_0 | v_601_0;
  assign v_2898_0 = v_607_0 | v_26_0;
  assign v_2899_0 = v_2900_0 | v_10685_0;
  assign v_2900_0 = v_2901_0 | v_10684_0;
  assign v_2901_0 = v_589_0 ? v_2902_0 : 3'h0;
  assign v_2903_0 = v_2904_0 | v_2905_0;
  assign v_2904_0 = v_589_0 | v_601_0;
  assign v_2905_0 = v_607_0 | v_26_0;
  assign v_2906_0 = v_2907_0 | v_10681_0;
  assign v_2907_0 = v_2908_0 | v_10680_0;
  assign v_2908_0 = v_589_0 ? v_2909_0 : 3'h0;
  assign v_2910_0 = v_2911_0 | v_2912_0;
  assign v_2911_0 = v_589_0 | v_601_0;
  assign v_2912_0 = v_607_0 | v_26_0;
  assign v_2913_0 = v_2914_0 | v_10677_0;
  assign v_2914_0 = v_2915_0 | v_10676_0;
  assign v_2915_0 = v_589_0 ? v_2916_0 : 3'h0;
  assign v_2917_0 = v_2918_0 | v_2919_0;
  assign v_2918_0 = v_589_0 | v_601_0;
  assign v_2919_0 = v_607_0 | v_26_0;
  assign v_2920_0 = v_2921_0 | v_10673_0;
  assign v_2921_0 = v_2922_0 | v_10672_0;
  assign v_2922_0 = v_589_0 ? v_2923_0 : 3'h0;
  assign v_2924_0 = v_2925_0 | v_2926_0;
  assign v_2925_0 = v_589_0 | v_601_0;
  assign v_2926_0 = v_607_0 | v_26_0;
  assign v_2927_0 = v_2928_0 | v_10669_0;
  assign v_2928_0 = v_2929_0 | v_10668_0;
  assign v_2929_0 = v_589_0 ? v_2930_0 : 3'h0;
  assign v_2931_0 = v_2932_0 | v_2933_0;
  assign v_2932_0 = v_589_0 | v_601_0;
  assign v_2933_0 = v_607_0 | v_26_0;
  assign v_2934_0 = v_2935_0 | v_10665_0;
  assign v_2935_0 = v_2936_0 | v_10664_0;
  assign v_2936_0 = v_589_0 ? v_2937_0 : 3'h0;
  assign v_2938_0 = v_2939_0 | v_2940_0;
  assign v_2939_0 = v_589_0 | v_601_0;
  assign v_2940_0 = v_607_0 | v_26_0;
  assign v_2941_0 = v_2942_0 | v_10661_0;
  assign v_2942_0 = v_2943_0 | v_10660_0;
  assign v_2943_0 = v_589_0 ? v_2944_0 : 3'h0;
  assign v_2945_0 = v_2946_0 | v_2947_0;
  assign v_2946_0 = v_589_0 | v_601_0;
  assign v_2947_0 = v_607_0 | v_26_0;
  assign v_2948_0 = v_2949_0 | v_10657_0;
  assign v_2949_0 = v_2950_0 | v_10656_0;
  assign v_2950_0 = v_589_0 ? v_2951_0 : 3'h0;
  assign v_2952_0 = v_2953_0 | v_2954_0;
  assign v_2953_0 = v_589_0 | v_601_0;
  assign v_2954_0 = v_607_0 | v_26_0;
  assign v_2955_0 = v_2956_0 | v_10653_0;
  assign v_2956_0 = v_2957_0 | v_10652_0;
  assign v_2957_0 = v_589_0 ? v_2958_0 : 3'h0;
  assign v_2959_0 = v_2960_0 | v_2961_0;
  assign v_2960_0 = v_589_0 | v_601_0;
  assign v_2961_0 = v_607_0 | v_26_0;
  assign v_2962_0 = v_2963_0 | v_10649_0;
  assign v_2963_0 = v_2964_0 | v_10648_0;
  assign v_2964_0 = v_589_0 ? v_2965_0 : 3'h0;
  assign v_2966_0 = v_2967_0 | v_2968_0;
  assign v_2967_0 = v_589_0 | v_601_0;
  assign v_2968_0 = v_607_0 | v_26_0;
  assign v_2969_0 = v_2970_0 | v_10645_0;
  assign v_2970_0 = v_2971_0 | v_10644_0;
  assign v_2971_0 = v_589_0 ? v_2972_0 : 3'h0;
  assign v_2973_0 = v_2974_0 | v_2975_0;
  assign v_2974_0 = v_589_0 | v_601_0;
  assign v_2975_0 = v_607_0 | v_26_0;
  assign v_2976_0 = v_2977_0 | v_10641_0;
  assign v_2977_0 = v_2978_0 | v_10640_0;
  assign v_2978_0 = v_589_0 ? v_2979_0 : 3'h0;
  assign v_2980_0 = v_2981_0 | v_2982_0;
  assign v_2981_0 = v_589_0 | v_601_0;
  assign v_2982_0 = v_607_0 | v_26_0;
  assign v_2983_0 = v_2984_0 | v_10637_0;
  assign v_2984_0 = v_2985_0 | v_10636_0;
  assign v_2985_0 = v_589_0 ? v_2986_0 : 3'h0;
  assign v_2987_0 = v_2988_0 | v_2989_0;
  assign v_2988_0 = v_589_0 | v_601_0;
  assign v_2989_0 = v_607_0 | v_26_0;
  assign v_2990_0 = v_2991_0 | v_10633_0;
  assign v_2991_0 = v_2992_0 | v_10632_0;
  assign v_2992_0 = v_589_0 ? v_2993_0 : 3'h0;
  assign v_2994_0 = v_2995_0 | v_2996_0;
  assign v_2995_0 = v_589_0 | v_601_0;
  assign v_2996_0 = v_607_0 | v_26_0;
  assign v_2997_0 = v_2998_0 | v_10629_0;
  assign v_2998_0 = v_2999_0 | v_10628_0;
  assign v_2999_0 = v_589_0 ? v_3000_0 : 3'h0;
  assign v_3001_0 = v_3002_0 | v_3003_0;
  assign v_3002_0 = v_589_0 | v_601_0;
  assign v_3003_0 = v_607_0 | v_26_0;
  assign v_3004_0 = v_3005_0 | v_10625_0;
  assign v_3005_0 = v_3006_0 | v_10624_0;
  assign v_3006_0 = v_589_0 ? v_3007_0 : 3'h0;
  assign v_3008_0 = v_3009_0 | v_3010_0;
  assign v_3009_0 = v_589_0 | v_601_0;
  assign v_3010_0 = v_607_0 | v_26_0;
  assign v_3011_0 = v_3012_0 | v_10621_0;
  assign v_3012_0 = v_3013_0 | v_10620_0;
  assign v_3013_0 = v_589_0 ? v_3014_0 : 3'h0;
  assign v_3015_0 = v_3016_0 | v_3017_0;
  assign v_3016_0 = v_589_0 | v_601_0;
  assign v_3017_0 = v_607_0 | v_26_0;
  assign v_3018_0 = v_3019_0 | v_10617_0;
  assign v_3019_0 = v_3020_0 | v_10616_0;
  assign v_3020_0 = v_589_0 ? v_3021_0 : 3'h0;
  assign v_3022_0 = v_3023_0 | v_3024_0;
  assign v_3023_0 = v_589_0 | v_601_0;
  assign v_3024_0 = v_607_0 | v_26_0;
  assign v_3025_0 = v_3026_0 | v_10613_0;
  assign v_3026_0 = v_3027_0 | v_10612_0;
  assign v_3027_0 = v_589_0 ? v_3028_0 : 3'h0;
  assign v_3029_0 = v_3030_0 | v_3031_0;
  assign v_3030_0 = v_589_0 | v_601_0;
  assign v_3031_0 = v_607_0 | v_26_0;
  assign v_3032_0 = v_3033_0 | v_10609_0;
  assign v_3033_0 = v_3034_0 | v_10608_0;
  assign v_3034_0 = v_589_0 ? v_3035_0 : 3'h0;
  assign v_3036_0 = v_3037_0 | v_3038_0;
  assign v_3037_0 = v_589_0 | v_601_0;
  assign v_3038_0 = v_607_0 | v_26_0;
  assign v_3039_0 = v_3040_0 | v_10605_0;
  assign v_3040_0 = v_3041_0 | v_10604_0;
  assign v_3041_0 = v_589_0 ? v_3042_0 : 3'h0;
  assign v_3043_0 = v_3044_0 | v_3045_0;
  assign v_3044_0 = v_589_0 | v_601_0;
  assign v_3045_0 = v_607_0 | v_26_0;
  assign v_3046_0 = v_3047_0 | v_10601_0;
  assign v_3047_0 = v_3048_0 | v_10600_0;
  assign v_3048_0 = v_589_0 ? v_3049_0 : 3'h0;
  assign v_3050_0 = v_3051_0 | v_3052_0;
  assign v_3051_0 = v_589_0 | v_601_0;
  assign v_3052_0 = v_607_0 | v_26_0;
  assign v_3053_0 = v_3054_0 | v_10597_0;
  assign v_3054_0 = v_3055_0 | v_10596_0;
  assign v_3055_0 = v_589_0 ? v_3056_0 : 3'h0;
  assign v_3057_0 = v_3058_0 | v_3059_0;
  assign v_3058_0 = v_589_0 | v_601_0;
  assign v_3059_0 = v_607_0 | v_26_0;
  assign v_3060_0 = v_3061_0 | v_10593_0;
  assign v_3061_0 = v_3062_0 | v_10592_0;
  assign v_3062_0 = v_589_0 ? v_3063_0 : 3'h0;
  assign v_3064_0 = v_3065_0 | v_3066_0;
  assign v_3065_0 = v_589_0 | v_601_0;
  assign v_3066_0 = v_607_0 | v_26_0;
  assign v_3067_0 = v_3068_0 | v_10589_0;
  assign v_3068_0 = v_3069_0 | v_10588_0;
  assign v_3069_0 = v_589_0 ? v_3070_0 : 3'h0;
  assign v_3071_0 = v_3072_0 | v_3073_0;
  assign v_3072_0 = v_589_0 | v_601_0;
  assign v_3073_0 = v_607_0 | v_26_0;
  assign v_3074_0 = v_3075_0 | v_10585_0;
  assign v_3075_0 = v_3076_0 | v_10584_0;
  assign v_3076_0 = v_589_0 ? v_3077_0 : 3'h0;
  assign v_3078_0 = v_3079_0 | v_3080_0;
  assign v_3079_0 = v_589_0 | v_601_0;
  assign v_3080_0 = v_607_0 | v_26_0;
  assign v_3081_0 = v_3082_0 | v_10581_0;
  assign v_3082_0 = v_3083_0 | v_10580_0;
  assign v_3083_0 = v_589_0 ? v_3084_0 : 3'h0;
  assign v_3085_0 = v_3086_0 | v_3087_0;
  assign v_3086_0 = v_589_0 | v_601_0;
  assign v_3087_0 = v_607_0 | v_26_0;
  assign v_3088_0 = v_3089_0 | v_10577_0;
  assign v_3089_0 = v_3090_0 | v_10576_0;
  assign v_3090_0 = v_589_0 ? v_3091_0 : 3'h0;
  assign v_3092_0 = v_3093_0 | v_3094_0;
  assign v_3093_0 = v_589_0 | v_601_0;
  assign v_3094_0 = v_607_0 | v_26_0;
  assign v_3095_0 = v_3096_0 | v_10573_0;
  assign v_3096_0 = v_3097_0 | v_10572_0;
  assign v_3097_0 = v_589_0 ? v_3098_0 : 3'h0;
  assign v_3099_0 = v_3100_0 | v_3101_0;
  assign v_3100_0 = v_589_0 | v_601_0;
  assign v_3101_0 = v_607_0 | v_26_0;
  assign v_3102_0 = v_3103_0 | v_10569_0;
  assign v_3103_0 = v_3104_0 | v_10568_0;
  assign v_3104_0 = v_589_0 ? v_3105_0 : 3'h0;
  assign v_3106_0 = v_3107_0 | v_3108_0;
  assign v_3107_0 = v_589_0 | v_601_0;
  assign v_3108_0 = v_607_0 | v_26_0;
  assign v_3109_0 = v_3110_0 | v_10565_0;
  assign v_3110_0 = v_3111_0 | v_10564_0;
  assign v_3111_0 = v_589_0 ? v_3112_0 : 3'h0;
  assign v_3113_0 = v_3114_0 | v_3115_0;
  assign v_3114_0 = v_589_0 | v_601_0;
  assign v_3115_0 = v_607_0 | v_26_0;
  assign v_3116_0 = v_3117_0 | v_10561_0;
  assign v_3117_0 = v_3118_0 | v_10560_0;
  assign v_3118_0 = v_589_0 ? v_3119_0 : 3'h0;
  assign v_3120_0 = v_3121_0 | v_3122_0;
  assign v_3121_0 = v_589_0 | v_601_0;
  assign v_3122_0 = v_607_0 | v_26_0;
  assign v_3123_0 = v_3124_0 | v_10557_0;
  assign v_3124_0 = v_3125_0 | v_10556_0;
  assign v_3125_0 = v_589_0 ? v_3126_0 : 3'h0;
  assign v_3127_0 = v_3128_0 | v_3129_0;
  assign v_3128_0 = v_589_0 | v_601_0;
  assign v_3129_0 = v_607_0 | v_26_0;
  assign v_3130_0 = v_3131_0 | v_10553_0;
  assign v_3131_0 = v_3132_0 | v_10552_0;
  assign v_3132_0 = v_589_0 ? v_3133_0 : 3'h0;
  assign v_3134_0 = v_3135_0 | v_3136_0;
  assign v_3135_0 = v_589_0 | v_601_0;
  assign v_3136_0 = v_607_0 | v_26_0;
  assign v_3137_0 = v_3138_0 | v_10549_0;
  assign v_3138_0 = v_3139_0 | v_10548_0;
  assign v_3139_0 = v_589_0 ? v_3140_0 : 3'h0;
  assign v_3141_0 = v_3142_0 | v_3143_0;
  assign v_3142_0 = v_589_0 | v_601_0;
  assign v_3143_0 = v_607_0 | v_26_0;
  assign v_3144_0 = v_3145_0 | v_10545_0;
  assign v_3145_0 = v_3146_0 | v_10544_0;
  assign v_3146_0 = v_589_0 ? v_3147_0 : 3'h0;
  assign v_3148_0 = v_3149_0 | v_3150_0;
  assign v_3149_0 = v_589_0 | v_601_0;
  assign v_3150_0 = v_607_0 | v_26_0;
  assign v_3151_0 = v_3152_0 | v_10541_0;
  assign v_3152_0 = v_3153_0 | v_10540_0;
  assign v_3153_0 = v_589_0 ? v_3154_0 : 3'h0;
  assign v_3155_0 = v_3156_0 | v_3157_0;
  assign v_3156_0 = v_589_0 | v_601_0;
  assign v_3157_0 = v_607_0 | v_26_0;
  assign v_3158_0 = v_3159_0 | v_10537_0;
  assign v_3159_0 = v_3160_0 | v_10536_0;
  assign v_3160_0 = v_589_0 ? v_3161_0 : 3'h0;
  assign v_3162_0 = v_3163_0 | v_3164_0;
  assign v_3163_0 = v_589_0 | v_601_0;
  assign v_3164_0 = v_607_0 | v_26_0;
  assign v_3165_0 = v_3166_0 | v_10533_0;
  assign v_3166_0 = v_3167_0 | v_10532_0;
  assign v_3167_0 = v_589_0 ? v_3168_0 : 3'h0;
  assign v_3169_0 = v_3170_0 | v_3171_0;
  assign v_3170_0 = v_589_0 | v_601_0;
  assign v_3171_0 = v_607_0 | v_26_0;
  assign v_3172_0 = v_3173_0 | v_10529_0;
  assign v_3173_0 = v_3174_0 | v_10528_0;
  assign v_3174_0 = v_589_0 ? v_3175_0 : 3'h0;
  assign v_3176_0 = v_3177_0 | v_3178_0;
  assign v_3177_0 = v_589_0 | v_601_0;
  assign v_3178_0 = v_607_0 | v_26_0;
  assign v_3179_0 = v_3180_0 | v_10525_0;
  assign v_3180_0 = v_3181_0 | v_10524_0;
  assign v_3181_0 = v_589_0 ? v_3182_0 : 3'h0;
  assign v_3183_0 = v_3184_0 | v_3185_0;
  assign v_3184_0 = v_589_0 | v_601_0;
  assign v_3185_0 = v_607_0 | v_26_0;
  assign v_3186_0 = v_3187_0 | v_10521_0;
  assign v_3187_0 = v_3188_0 | v_10520_0;
  assign v_3188_0 = v_589_0 ? v_3189_0 : 3'h0;
  assign v_3190_0 = v_3191_0 | v_3192_0;
  assign v_3191_0 = v_589_0 | v_601_0;
  assign v_3192_0 = v_607_0 | v_26_0;
  assign v_3193_0 = v_3194_0 | v_10517_0;
  assign v_3194_0 = v_3195_0 | v_10516_0;
  assign v_3195_0 = v_589_0 ? v_3196_0 : 3'h0;
  assign v_3197_0 = v_3198_0 | v_3199_0;
  assign v_3198_0 = v_589_0 | v_601_0;
  assign v_3199_0 = v_607_0 | v_26_0;
  assign v_3200_0 = v_3201_0 | v_10513_0;
  assign v_3201_0 = v_3202_0 | v_10512_0;
  assign v_3202_0 = v_589_0 ? v_3203_0 : 3'h0;
  assign v_3204_0 = v_3205_0 | v_3206_0;
  assign v_3205_0 = v_589_0 | v_601_0;
  assign v_3206_0 = v_607_0 | v_26_0;
  assign v_3207_0 = v_3208_0 | v_10509_0;
  assign v_3208_0 = v_3209_0 | v_10508_0;
  assign v_3209_0 = v_589_0 ? v_3210_0 : 3'h0;
  assign v_3211_0 = v_3212_0 | v_3213_0;
  assign v_3212_0 = v_589_0 | v_601_0;
  assign v_3213_0 = v_607_0 | v_26_0;
  assign v_3214_0 = v_3215_0 | v_10505_0;
  assign v_3215_0 = v_3216_0 | v_10504_0;
  assign v_3216_0 = v_589_0 ? v_3217_0 : 3'h0;
  assign v_3218_0 = v_3219_0 | v_3220_0;
  assign v_3219_0 = v_589_0 | v_601_0;
  assign v_3220_0 = v_607_0 | v_26_0;
  assign v_3221_0 = v_3222_0 | v_10501_0;
  assign v_3222_0 = v_3223_0 | v_10500_0;
  assign v_3223_0 = v_589_0 ? v_3224_0 : 3'h0;
  assign v_3225_0 = v_3226_0 | v_3227_0;
  assign v_3226_0 = v_589_0 | v_601_0;
  assign v_3227_0 = v_607_0 | v_26_0;
  assign v_3228_0 = v_3229_0 | v_10497_0;
  assign v_3229_0 = v_3230_0 | v_10496_0;
  assign v_3230_0 = v_589_0 ? v_3231_0 : 3'h0;
  assign v_3232_0 = v_3233_0 | v_3234_0;
  assign v_3233_0 = v_589_0 | v_601_0;
  assign v_3234_0 = v_607_0 | v_26_0;
  assign v_3235_0 = v_3236_0 | v_10493_0;
  assign v_3236_0 = v_3237_0 | v_10492_0;
  assign v_3237_0 = v_589_0 ? v_3238_0 : 3'h0;
  assign v_3239_0 = v_3240_0 | v_3241_0;
  assign v_3240_0 = v_589_0 | v_601_0;
  assign v_3241_0 = v_607_0 | v_26_0;
  assign v_3242_0 = v_3243_0 | v_10489_0;
  assign v_3243_0 = v_3244_0 | v_10488_0;
  assign v_3244_0 = v_589_0 ? v_3245_0 : 3'h0;
  assign v_3246_0 = v_3247_0 | v_3248_0;
  assign v_3247_0 = v_589_0 | v_601_0;
  assign v_3248_0 = v_607_0 | v_26_0;
  assign v_3249_0 = v_3250_0 | v_10485_0;
  assign v_3250_0 = v_3251_0 | v_10484_0;
  assign v_3251_0 = v_589_0 ? v_3252_0 : 3'h0;
  assign v_3253_0 = v_3254_0 | v_3255_0;
  assign v_3254_0 = v_589_0 | v_601_0;
  assign v_3255_0 = v_607_0 | v_26_0;
  assign v_3256_0 = v_3257_0 | v_10481_0;
  assign v_3257_0 = v_3258_0 | v_10480_0;
  assign v_3258_0 = v_589_0 ? v_3259_0 : 3'h0;
  assign v_3260_0 = v_3261_0 | v_3262_0;
  assign v_3261_0 = v_589_0 | v_601_0;
  assign v_3262_0 = v_607_0 | v_26_0;
  assign v_3263_0 = v_3264_0 | v_10477_0;
  assign v_3264_0 = v_3265_0 | v_10476_0;
  assign v_3265_0 = v_589_0 ? v_3266_0 : 3'h0;
  assign v_3267_0 = v_3268_0 | v_3269_0;
  assign v_3268_0 = v_589_0 | v_601_0;
  assign v_3269_0 = v_607_0 | v_26_0;
  assign v_3270_0 = v_3271_0 | v_10473_0;
  assign v_3271_0 = v_3272_0 | v_10472_0;
  assign v_3272_0 = v_589_0 ? v_3273_0 : 3'h0;
  assign v_3274_0 = v_3275_0 | v_3276_0;
  assign v_3275_0 = v_589_0 | v_601_0;
  assign v_3276_0 = v_607_0 | v_26_0;
  assign v_3277_0 = v_3278_0 | v_10469_0;
  assign v_3278_0 = v_3279_0 | v_10468_0;
  assign v_3279_0 = v_589_0 ? v_3280_0 : 3'h0;
  assign v_3281_0 = v_3282_0 | v_3283_0;
  assign v_3282_0 = v_589_0 | v_601_0;
  assign v_3283_0 = v_607_0 | v_26_0;
  assign v_3284_0 = v_3285_0 | v_10465_0;
  assign v_3285_0 = v_3286_0 | v_10464_0;
  assign v_3286_0 = v_589_0 ? v_3287_0 : 3'h0;
  assign v_3288_0 = v_3289_0 | v_3290_0;
  assign v_3289_0 = v_589_0 | v_601_0;
  assign v_3290_0 = v_607_0 | v_26_0;
  assign v_3291_0 = v_3292_0 | v_10461_0;
  assign v_3292_0 = v_3293_0 | v_10460_0;
  assign v_3293_0 = v_589_0 ? v_3294_0 : 3'h0;
  assign v_3295_0 = v_3296_0 | v_3297_0;
  assign v_3296_0 = v_589_0 | v_601_0;
  assign v_3297_0 = v_607_0 | v_26_0;
  assign v_3298_0 = v_3299_0 | v_10457_0;
  assign v_3299_0 = v_3300_0 | v_10456_0;
  assign v_3300_0 = v_589_0 ? v_3301_0 : 3'h0;
  assign v_3302_0 = v_3303_0 | v_3304_0;
  assign v_3303_0 = v_589_0 | v_601_0;
  assign v_3304_0 = v_607_0 | v_26_0;
  assign v_3305_0 = v_3306_0 | v_10453_0;
  assign v_3306_0 = v_3307_0 | v_10452_0;
  assign v_3307_0 = v_589_0 ? v_3308_0 : 3'h0;
  assign v_3309_0 = v_3310_0 | v_3311_0;
  assign v_3310_0 = v_589_0 | v_601_0;
  assign v_3311_0 = v_607_0 | v_26_0;
  assign v_3312_0 = v_3313_0 | v_10449_0;
  assign v_3313_0 = v_3314_0 | v_10448_0;
  assign v_3314_0 = v_589_0 ? v_3315_0 : 3'h0;
  assign v_3316_0 = v_3317_0 | v_3318_0;
  assign v_3317_0 = v_589_0 | v_601_0;
  assign v_3318_0 = v_607_0 | v_26_0;
  assign v_3319_0 = v_3320_0 | v_10445_0;
  assign v_3320_0 = v_3321_0 | v_10444_0;
  assign v_3321_0 = v_589_0 ? v_3322_0 : 3'h0;
  assign v_3323_0 = v_3324_0 | v_3325_0;
  assign v_3324_0 = v_589_0 | v_601_0;
  assign v_3325_0 = v_607_0 | v_26_0;
  assign v_3326_0 = v_3327_0 | v_10441_0;
  assign v_3327_0 = v_3328_0 | v_10440_0;
  assign v_3328_0 = v_589_0 ? v_3329_0 : 3'h0;
  assign v_3330_0 = v_3331_0 | v_3332_0;
  assign v_3331_0 = v_589_0 | v_601_0;
  assign v_3332_0 = v_607_0 | v_26_0;
  assign v_3333_0 = v_3334_0 | v_10437_0;
  assign v_3334_0 = v_3335_0 | v_10436_0;
  assign v_3335_0 = v_589_0 ? v_3336_0 : 3'h0;
  assign v_3337_0 = v_3338_0 | v_3339_0;
  assign v_3338_0 = v_589_0 | v_601_0;
  assign v_3339_0 = v_607_0 | v_26_0;
  assign v_3340_0 = v_3341_0 | v_10433_0;
  assign v_3341_0 = v_3342_0 | v_10432_0;
  assign v_3342_0 = v_589_0 ? v_3343_0 : 3'h0;
  assign v_3344_0 = v_3345_0 | v_3346_0;
  assign v_3345_0 = v_589_0 | v_601_0;
  assign v_3346_0 = v_607_0 | v_26_0;
  assign v_3347_0 = v_3348_0 | v_10429_0;
  assign v_3348_0 = v_3349_0 | v_10428_0;
  assign v_3349_0 = v_589_0 ? v_3350_0 : 3'h0;
  assign v_3351_0 = v_3352_0 | v_3353_0;
  assign v_3352_0 = v_589_0 | v_601_0;
  assign v_3353_0 = v_607_0 | v_26_0;
  assign v_3354_0 = v_3355_0 | v_10425_0;
  assign v_3355_0 = v_3356_0 | v_10424_0;
  assign v_3356_0 = v_589_0 ? v_3357_0 : 3'h0;
  assign v_3358_0 = v_3359_0 | v_3360_0;
  assign v_3359_0 = v_589_0 | v_601_0;
  assign v_3360_0 = v_607_0 | v_26_0;
  assign v_3361_0 = v_3362_0 | v_10421_0;
  assign v_3362_0 = v_3363_0 | v_10420_0;
  assign v_3363_0 = v_589_0 ? v_3364_0 : 3'h0;
  assign v_3365_0 = v_3366_0 | v_3367_0;
  assign v_3366_0 = v_589_0 | v_601_0;
  assign v_3367_0 = v_607_0 | v_26_0;
  assign v_3368_0 = v_3369_0 | v_10417_0;
  assign v_3369_0 = v_3370_0 | v_10416_0;
  assign v_3370_0 = v_589_0 ? v_3371_0 : 3'h0;
  assign v_3372_0 = v_3373_0 | v_3374_0;
  assign v_3373_0 = v_589_0 | v_601_0;
  assign v_3374_0 = v_607_0 | v_26_0;
  assign v_3375_0 = v_3376_0 | v_10413_0;
  assign v_3376_0 = v_3377_0 | v_10412_0;
  assign v_3377_0 = v_589_0 ? v_3378_0 : 3'h0;
  assign v_3379_0 = v_3380_0 | v_3381_0;
  assign v_3380_0 = v_589_0 | v_601_0;
  assign v_3381_0 = v_607_0 | v_26_0;
  assign v_3382_0 = v_3383_0 | v_10409_0;
  assign v_3383_0 = v_3384_0 | v_10408_0;
  assign v_3384_0 = v_589_0 ? v_3385_0 : 3'h0;
  assign v_3386_0 = v_3387_0 | v_3388_0;
  assign v_3387_0 = v_589_0 | v_601_0;
  assign v_3388_0 = v_607_0 | v_26_0;
  assign v_3389_0 = v_3390_0 | v_10405_0;
  assign v_3390_0 = v_3391_0 | v_10404_0;
  assign v_3391_0 = v_589_0 ? v_3392_0 : 3'h0;
  assign v_3393_0 = v_3394_0 | v_3395_0;
  assign v_3394_0 = v_589_0 | v_601_0;
  assign v_3395_0 = v_607_0 | v_26_0;
  assign v_3396_0 = v_3397_0 | v_10401_0;
  assign v_3397_0 = v_3398_0 | v_10400_0;
  assign v_3398_0 = v_589_0 ? v_3399_0 : 3'h0;
  assign v_3400_0 = v_3401_0 | v_3402_0;
  assign v_3401_0 = v_589_0 | v_601_0;
  assign v_3402_0 = v_607_0 | v_26_0;
  assign v_3403_0 = v_3404_0 | v_10397_0;
  assign v_3404_0 = v_3405_0 | v_10396_0;
  assign v_3405_0 = v_589_0 ? v_3406_0 : 3'h0;
  assign v_3407_0 = v_3408_0 | v_3409_0;
  assign v_3408_0 = v_589_0 | v_601_0;
  assign v_3409_0 = v_607_0 | v_26_0;
  assign v_3410_0 = v_3411_0 | v_10393_0;
  assign v_3411_0 = v_3412_0 | v_10392_0;
  assign v_3412_0 = v_589_0 ? v_3413_0 : 3'h0;
  assign v_3414_0 = v_3415_0 | v_3416_0;
  assign v_3415_0 = v_589_0 | v_601_0;
  assign v_3416_0 = v_607_0 | v_26_0;
  assign v_3417_0 = v_3418_0 | v_10389_0;
  assign v_3418_0 = v_3419_0 | v_10388_0;
  assign v_3419_0 = v_589_0 ? v_3420_0 : 3'h0;
  assign v_3421_0 = v_3422_0 | v_3423_0;
  assign v_3422_0 = v_589_0 | v_601_0;
  assign v_3423_0 = v_607_0 | v_26_0;
  assign v_3424_0 = v_3425_0 | v_10385_0;
  assign v_3425_0 = v_3426_0 | v_10384_0;
  assign v_3426_0 = v_589_0 ? v_3427_0 : 3'h0;
  assign v_3428_0 = v_3429_0 | v_3430_0;
  assign v_3429_0 = v_589_0 | v_601_0;
  assign v_3430_0 = v_607_0 | v_26_0;
  assign v_3431_0 = v_3432_0 | v_10381_0;
  assign v_3432_0 = v_3433_0 | v_10380_0;
  assign v_3433_0 = v_589_0 ? v_3434_0 : 3'h0;
  assign v_3435_0 = v_3436_0 | v_3437_0;
  assign v_3436_0 = v_589_0 | v_601_0;
  assign v_3437_0 = v_607_0 | v_26_0;
  assign v_3438_0 = v_3439_0 | v_10377_0;
  assign v_3439_0 = v_3440_0 | v_10376_0;
  assign v_3440_0 = v_589_0 ? v_3441_0 : 3'h0;
  assign v_3442_0 = v_3443_0 | v_3444_0;
  assign v_3443_0 = v_589_0 | v_601_0;
  assign v_3444_0 = v_607_0 | v_26_0;
  assign v_3445_0 = v_3446_0 | v_10373_0;
  assign v_3446_0 = v_3447_0 | v_10372_0;
  assign v_3447_0 = v_589_0 ? v_3448_0 : 3'h0;
  assign v_3449_0 = v_3450_0 | v_3451_0;
  assign v_3450_0 = v_589_0 | v_601_0;
  assign v_3451_0 = v_607_0 | v_26_0;
  assign v_3452_0 = v_3453_0 | v_10369_0;
  assign v_3453_0 = v_3454_0 | v_10368_0;
  assign v_3454_0 = v_589_0 ? v_3455_0 : 3'h0;
  assign v_3456_0 = v_3457_0 | v_3458_0;
  assign v_3457_0 = v_589_0 | v_601_0;
  assign v_3458_0 = v_607_0 | v_26_0;
  assign v_3459_0 = v_3460_0 | v_10365_0;
  assign v_3460_0 = v_3461_0 | v_10364_0;
  assign v_3461_0 = v_589_0 ? v_3462_0 : 3'h0;
  assign v_3463_0 = v_3464_0 | v_3465_0;
  assign v_3464_0 = v_589_0 | v_601_0;
  assign v_3465_0 = v_607_0 | v_26_0;
  assign v_3466_0 = v_3467_0 | v_10361_0;
  assign v_3467_0 = v_3468_0 | v_10360_0;
  assign v_3468_0 = v_589_0 ? v_3469_0 : 3'h0;
  assign v_3470_0 = v_3471_0 | v_3472_0;
  assign v_3471_0 = v_589_0 | v_601_0;
  assign v_3472_0 = v_607_0 | v_26_0;
  assign v_3473_0 = v_3474_0 | v_10357_0;
  assign v_3474_0 = v_3475_0 | v_10356_0;
  assign v_3475_0 = v_589_0 ? v_3476_0 : 3'h0;
  assign v_3477_0 = v_3478_0 | v_3479_0;
  assign v_3478_0 = v_589_0 | v_601_0;
  assign v_3479_0 = v_607_0 | v_26_0;
  assign v_3480_0 = v_3481_0 | v_10353_0;
  assign v_3481_0 = v_3482_0 | v_10352_0;
  assign v_3482_0 = v_589_0 ? v_3483_0 : 3'h0;
  assign v_3484_0 = v_3485_0 | v_3486_0;
  assign v_3485_0 = v_589_0 | v_601_0;
  assign v_3486_0 = v_607_0 | v_26_0;
  assign v_3487_0 = v_3488_0 | v_10349_0;
  assign v_3488_0 = v_3489_0 | v_10348_0;
  assign v_3489_0 = v_589_0 ? v_3490_0 : 3'h0;
  assign v_3491_0 = v_3492_0 | v_3493_0;
  assign v_3492_0 = v_589_0 | v_601_0;
  assign v_3493_0 = v_607_0 | v_26_0;
  assign v_3494_0 = v_3495_0 | v_10345_0;
  assign v_3495_0 = v_3496_0 | v_10344_0;
  assign v_3496_0 = v_589_0 ? v_3497_0 : 3'h0;
  assign v_3498_0 = v_3499_0 | v_3500_0;
  assign v_3499_0 = v_589_0 | v_601_0;
  assign v_3500_0 = v_607_0 | v_26_0;
  assign v_3501_0 = v_3502_0 | v_10341_0;
  assign v_3502_0 = v_3503_0 | v_10340_0;
  assign v_3503_0 = v_589_0 ? v_3504_0 : 3'h0;
  assign v_3505_0 = v_3506_0 | v_3507_0;
  assign v_3506_0 = v_589_0 | v_601_0;
  assign v_3507_0 = v_607_0 | v_26_0;
  assign v_3508_0 = v_3509_0 | v_10337_0;
  assign v_3509_0 = v_3510_0 | v_10336_0;
  assign v_3510_0 = v_589_0 ? v_3511_0 : 3'h0;
  assign v_3512_0 = v_3513_0 | v_3514_0;
  assign v_3513_0 = v_589_0 | v_601_0;
  assign v_3514_0 = v_607_0 | v_26_0;
  assign v_3515_0 = v_3516_0 | v_10333_0;
  assign v_3516_0 = v_3517_0 | v_10332_0;
  assign v_3517_0 = v_589_0 ? v_3518_0 : 3'h0;
  assign v_3519_0 = v_3520_0 | v_3521_0;
  assign v_3520_0 = v_589_0 | v_601_0;
  assign v_3521_0 = v_607_0 | v_26_0;
  assign v_3522_0 = v_3523_0 | v_10329_0;
  assign v_3523_0 = v_3524_0 | v_10328_0;
  assign v_3524_0 = v_589_0 ? v_3525_0 : 3'h0;
  assign v_3526_0 = v_3527_0 | v_3528_0;
  assign v_3527_0 = v_589_0 | v_601_0;
  assign v_3528_0 = v_607_0 | v_26_0;
  assign v_3529_0 = v_3530_0 | v_10325_0;
  assign v_3530_0 = v_3531_0 | v_10324_0;
  assign v_3531_0 = v_589_0 ? v_3532_0 : 3'h0;
  assign v_3533_0 = v_3534_0 | v_3535_0;
  assign v_3534_0 = v_589_0 | v_601_0;
  assign v_3535_0 = v_607_0 | v_26_0;
  assign v_3536_0 = v_3537_0 | v_10321_0;
  assign v_3537_0 = v_3538_0 | v_10320_0;
  assign v_3538_0 = v_589_0 ? v_3539_0 : 3'h0;
  assign v_3540_0 = v_3541_0 | v_3542_0;
  assign v_3541_0 = v_589_0 | v_601_0;
  assign v_3542_0 = v_607_0 | v_26_0;
  assign v_3543_0 = v_3544_0 | v_10317_0;
  assign v_3544_0 = v_3545_0 | v_10316_0;
  assign v_3545_0 = v_589_0 ? v_3546_0 : 3'h0;
  assign v_3547_0 = v_3548_0 | v_3549_0;
  assign v_3548_0 = v_589_0 | v_601_0;
  assign v_3549_0 = v_607_0 | v_26_0;
  assign v_3550_0 = v_3551_0 | v_10313_0;
  assign v_3551_0 = v_3552_0 | v_10312_0;
  assign v_3552_0 = v_589_0 ? v_3553_0 : 3'h0;
  assign v_3554_0 = v_3555_0 | v_3556_0;
  assign v_3555_0 = v_589_0 | v_601_0;
  assign v_3556_0 = v_607_0 | v_26_0;
  assign v_3557_0 = v_3558_0 | v_10309_0;
  assign v_3558_0 = v_3559_0 | v_10308_0;
  assign v_3559_0 = v_589_0 ? v_3560_0 : 3'h0;
  assign v_3561_0 = v_3562_0 | v_3563_0;
  assign v_3562_0 = v_589_0 | v_601_0;
  assign v_3563_0 = v_607_0 | v_26_0;
  assign v_3564_0 = v_3565_0 | v_10305_0;
  assign v_3565_0 = v_3566_0 | v_10304_0;
  assign v_3566_0 = v_589_0 ? v_3567_0 : 3'h0;
  assign v_3568_0 = v_3569_0 | v_3570_0;
  assign v_3569_0 = v_589_0 | v_601_0;
  assign v_3570_0 = v_607_0 | v_26_0;
  assign v_3571_0 = v_3572_0 | v_10301_0;
  assign v_3572_0 = v_3573_0 | v_10300_0;
  assign v_3573_0 = v_589_0 ? v_3574_0 : 3'h0;
  assign v_3575_0 = v_3576_0 | v_3577_0;
  assign v_3576_0 = v_589_0 | v_601_0;
  assign v_3577_0 = v_607_0 | v_26_0;
  assign v_3578_0 = v_3579_0 | v_10297_0;
  assign v_3579_0 = v_3580_0 | v_10296_0;
  assign v_3580_0 = v_589_0 ? v_3581_0 : 3'h0;
  assign v_3582_0 = v_3583_0 | v_3584_0;
  assign v_3583_0 = v_589_0 | v_601_0;
  assign v_3584_0 = v_607_0 | v_26_0;
  assign v_3585_0 = v_3586_0 | v_10293_0;
  assign v_3586_0 = v_3587_0 | v_10292_0;
  assign v_3587_0 = v_589_0 ? v_3588_0 : 3'h0;
  assign v_3589_0 = v_3590_0 | v_3591_0;
  assign v_3590_0 = v_589_0 | v_601_0;
  assign v_3591_0 = v_607_0 | v_26_0;
  assign v_3592_0 = v_3593_0 | v_10289_0;
  assign v_3593_0 = v_3594_0 | v_10288_0;
  assign v_3594_0 = v_589_0 ? v_3595_0 : 3'h0;
  assign v_3596_0 = v_3597_0 | v_3598_0;
  assign v_3597_0 = v_589_0 | v_601_0;
  assign v_3598_0 = v_607_0 | v_26_0;
  assign v_3599_0 = v_3600_0 | v_10285_0;
  assign v_3600_0 = v_3601_0 | v_10284_0;
  assign v_3601_0 = v_589_0 ? v_3602_0 : 3'h0;
  assign v_3603_0 = v_3604_0 | v_3605_0;
  assign v_3604_0 = v_589_0 | v_601_0;
  assign v_3605_0 = v_607_0 | v_26_0;
  assign v_3606_0 = v_3607_0 | v_10281_0;
  assign v_3607_0 = v_3608_0 | v_10280_0;
  assign v_3608_0 = v_589_0 ? v_3609_0 : 3'h0;
  assign v_3610_0 = v_3611_0 | v_3612_0;
  assign v_3611_0 = v_589_0 | v_601_0;
  assign v_3612_0 = v_607_0 | v_26_0;
  assign v_3613_0 = v_3614_0 | v_10277_0;
  assign v_3614_0 = v_3615_0 | v_10276_0;
  assign v_3615_0 = v_589_0 ? v_3616_0 : 3'h0;
  assign v_3617_0 = v_3618_0 | v_3619_0;
  assign v_3618_0 = v_589_0 | v_601_0;
  assign v_3619_0 = v_607_0 | v_26_0;
  assign v_3620_0 = v_3621_0 | v_10273_0;
  assign v_3621_0 = v_3622_0 | v_10272_0;
  assign v_3622_0 = v_589_0 ? v_3623_0 : 3'h0;
  assign v_3624_0 = v_3625_0 | v_3626_0;
  assign v_3625_0 = v_589_0 | v_601_0;
  assign v_3626_0 = v_607_0 | v_26_0;
  assign v_3627_0 = v_3628_0 | v_10269_0;
  assign v_3628_0 = v_3629_0 | v_10268_0;
  assign v_3629_0 = v_589_0 ? v_3630_0 : 3'h0;
  assign v_3631_0 = v_3632_0 | v_3633_0;
  assign v_3632_0 = v_589_0 | v_601_0;
  assign v_3633_0 = v_607_0 | v_26_0;
  assign v_3634_0 = v_3635_0 | v_10265_0;
  assign v_3635_0 = v_3636_0 | v_10264_0;
  assign v_3636_0 = v_589_0 ? v_3637_0 : 3'h0;
  assign v_3638_0 = v_3639_0 | v_3640_0;
  assign v_3639_0 = v_589_0 | v_601_0;
  assign v_3640_0 = v_607_0 | v_26_0;
  assign v_3641_0 = v_3642_0 | v_10261_0;
  assign v_3642_0 = v_3643_0 | v_10260_0;
  assign v_3643_0 = v_589_0 ? v_3644_0 : 3'h0;
  assign v_3645_0 = v_3646_0 | v_3647_0;
  assign v_3646_0 = v_589_0 | v_601_0;
  assign v_3647_0 = v_607_0 | v_26_0;
  assign v_3648_0 = v_3649_0 | v_10257_0;
  assign v_3649_0 = v_3650_0 | v_10256_0;
  assign v_3650_0 = v_589_0 ? v_3651_0 : 3'h0;
  assign v_3652_0 = v_3653_0 | v_3654_0;
  assign v_3653_0 = v_589_0 | v_601_0;
  assign v_3654_0 = v_607_0 | v_26_0;
  assign v_3655_0 = v_3656_0 | v_10253_0;
  assign v_3656_0 = v_3657_0 | v_10252_0;
  assign v_3657_0 = v_589_0 ? v_3658_0 : 3'h0;
  assign v_3659_0 = v_3660_0 | v_3661_0;
  assign v_3660_0 = v_589_0 | v_601_0;
  assign v_3661_0 = v_607_0 | v_26_0;
  assign v_3662_0 = v_3663_0 | v_10249_0;
  assign v_3663_0 = v_3664_0 | v_10248_0;
  assign v_3664_0 = v_589_0 ? v_3665_0 : 3'h0;
  assign v_3666_0 = v_3667_0 | v_3668_0;
  assign v_3667_0 = v_589_0 | v_601_0;
  assign v_3668_0 = v_607_0 | v_26_0;
  assign v_3669_0 = v_3670_0 | v_10245_0;
  assign v_3670_0 = v_3671_0 | v_10244_0;
  assign v_3671_0 = v_589_0 ? v_3672_0 : 3'h0;
  assign v_3673_0 = v_3674_0 | v_3675_0;
  assign v_3674_0 = v_589_0 | v_601_0;
  assign v_3675_0 = v_607_0 | v_26_0;
  assign v_3676_0 = v_3677_0 | v_10241_0;
  assign v_3677_0 = v_3678_0 | v_10240_0;
  assign v_3678_0 = v_589_0 ? v_3679_0 : 3'h0;
  assign v_3680_0 = v_3681_0 | v_3682_0;
  assign v_3681_0 = v_589_0 | v_601_0;
  assign v_3682_0 = v_607_0 | v_26_0;
  assign v_3683_0 = v_3684_0 | v_10237_0;
  assign v_3684_0 = v_3685_0 | v_10236_0;
  assign v_3685_0 = v_589_0 ? v_3686_0 : 3'h0;
  assign v_3687_0 = v_3688_0 | v_3689_0;
  assign v_3688_0 = v_589_0 | v_601_0;
  assign v_3689_0 = v_607_0 | v_26_0;
  assign v_3690_0 = v_3691_0 | v_10233_0;
  assign v_3691_0 = v_3692_0 | v_10232_0;
  assign v_3692_0 = v_589_0 ? v_3693_0 : 3'h0;
  assign v_3694_0 = v_3695_0 | v_3696_0;
  assign v_3695_0 = v_589_0 | v_601_0;
  assign v_3696_0 = v_607_0 | v_26_0;
  assign v_3697_0 = v_3698_0 | v_10229_0;
  assign v_3698_0 = v_3699_0 | v_10228_0;
  assign v_3699_0 = v_589_0 ? v_3700_0 : 3'h0;
  assign v_3701_0 = v_3702_0 | v_3703_0;
  assign v_3702_0 = v_589_0 | v_601_0;
  assign v_3703_0 = v_607_0 | v_26_0;
  assign v_3704_0 = v_3705_0 | v_10225_0;
  assign v_3705_0 = v_3706_0 | v_10224_0;
  assign v_3706_0 = v_589_0 ? v_3707_0 : 3'h0;
  assign v_3708_0 = v_3709_0 | v_3710_0;
  assign v_3709_0 = v_589_0 | v_601_0;
  assign v_3710_0 = v_607_0 | v_26_0;
  assign v_3711_0 = v_3712_0 | v_10221_0;
  assign v_3712_0 = v_3713_0 | v_10220_0;
  assign v_3713_0 = v_589_0 ? v_3714_0 : 3'h0;
  assign v_3715_0 = v_3716_0 | v_3717_0;
  assign v_3716_0 = v_589_0 | v_601_0;
  assign v_3717_0 = v_607_0 | v_26_0;
  assign v_3718_0 = v_3719_0 | v_10217_0;
  assign v_3719_0 = v_3720_0 | v_10216_0;
  assign v_3720_0 = v_589_0 ? v_3721_0 : 3'h0;
  assign v_3722_0 = v_3723_0 | v_3724_0;
  assign v_3723_0 = v_589_0 | v_601_0;
  assign v_3724_0 = v_607_0 | v_26_0;
  assign v_3725_0 = v_3726_0 | v_10213_0;
  assign v_3726_0 = v_3727_0 | v_10212_0;
  assign v_3727_0 = v_589_0 ? v_3728_0 : 3'h0;
  assign v_3729_0 = v_3730_0 | v_3731_0;
  assign v_3730_0 = v_589_0 | v_601_0;
  assign v_3731_0 = v_607_0 | v_26_0;
  assign v_3732_0 = v_3733_0 | v_10209_0;
  assign v_3733_0 = v_3734_0 | v_10208_0;
  assign v_3734_0 = v_589_0 ? v_3735_0 : 3'h0;
  assign v_3736_0 = v_3737_0 | v_3738_0;
  assign v_3737_0 = v_589_0 | v_601_0;
  assign v_3738_0 = v_607_0 | v_26_0;
  assign v_3739_0 = v_3740_0 | v_10205_0;
  assign v_3740_0 = v_3741_0 | v_10204_0;
  assign v_3741_0 = v_589_0 ? v_3742_0 : 3'h0;
  assign v_3743_0 = v_3744_0 | v_3745_0;
  assign v_3744_0 = v_589_0 | v_601_0;
  assign v_3745_0 = v_607_0 | v_26_0;
  assign v_3746_0 = v_3747_0 | v_10201_0;
  assign v_3747_0 = v_3748_0 | v_10200_0;
  assign v_3748_0 = v_589_0 ? v_3749_0 : 3'h0;
  assign v_3750_0 = v_3751_0 | v_3752_0;
  assign v_3751_0 = v_589_0 | v_601_0;
  assign v_3752_0 = v_607_0 | v_26_0;
  assign v_3753_0 = v_3754_0 | v_10197_0;
  assign v_3754_0 = v_3755_0 | v_10196_0;
  assign v_3755_0 = v_589_0 ? v_3756_0 : 3'h0;
  assign v_3757_0 = v_3758_0 | v_3759_0;
  assign v_3758_0 = v_589_0 | v_601_0;
  assign v_3759_0 = v_607_0 | v_26_0;
  assign v_3760_0 = v_3761_0 | v_10193_0;
  assign v_3761_0 = v_3762_0 | v_10192_0;
  assign v_3762_0 = v_589_0 ? v_3763_0 : 3'h0;
  assign v_3764_0 = v_3765_0 | v_3766_0;
  assign v_3765_0 = v_589_0 | v_601_0;
  assign v_3766_0 = v_607_0 | v_26_0;
  assign v_3767_0 = v_3768_0 | v_10189_0;
  assign v_3768_0 = v_3769_0 | v_10188_0;
  assign v_3769_0 = v_589_0 ? v_3770_0 : 3'h0;
  assign v_3771_0 = v_3772_0 | v_3773_0;
  assign v_3772_0 = v_589_0 | v_601_0;
  assign v_3773_0 = v_607_0 | v_26_0;
  assign v_3774_0 = v_3775_0 | v_10185_0;
  assign v_3775_0 = v_3776_0 | v_10184_0;
  assign v_3776_0 = v_589_0 ? v_3777_0 : 3'h0;
  assign v_3778_0 = v_3779_0 | v_3780_0;
  assign v_3779_0 = v_589_0 | v_601_0;
  assign v_3780_0 = v_607_0 | v_26_0;
  assign v_3781_0 = v_3782_0 | v_10181_0;
  assign v_3782_0 = v_3783_0 | v_10180_0;
  assign v_3783_0 = v_589_0 ? v_3784_0 : 3'h0;
  assign v_3785_0 = v_3786_0 | v_3787_0;
  assign v_3786_0 = v_589_0 | v_601_0;
  assign v_3787_0 = v_607_0 | v_26_0;
  assign v_3788_0 = v_3789_0 | v_10177_0;
  assign v_3789_0 = v_3790_0 | v_10176_0;
  assign v_3790_0 = v_589_0 ? v_3791_0 : 3'h0;
  assign v_3792_0 = v_3793_0 | v_3794_0;
  assign v_3793_0 = v_589_0 | v_601_0;
  assign v_3794_0 = v_607_0 | v_26_0;
  assign v_3795_0 = v_3796_0 | v_10173_0;
  assign v_3796_0 = v_3797_0 | v_10172_0;
  assign v_3797_0 = v_589_0 ? v_3798_0 : 3'h0;
  assign v_3799_0 = v_3800_0 | v_3801_0;
  assign v_3800_0 = v_589_0 | v_601_0;
  assign v_3801_0 = v_607_0 | v_26_0;
  assign v_3802_0 = v_3803_0 | v_10169_0;
  assign v_3803_0 = v_3804_0 | v_10168_0;
  assign v_3804_0 = v_589_0 ? v_3805_0 : 3'h0;
  assign v_3806_0 = v_3807_0 | v_3808_0;
  assign v_3807_0 = v_589_0 | v_601_0;
  assign v_3808_0 = v_607_0 | v_26_0;
  assign v_3809_0 = v_3810_0 | v_10165_0;
  assign v_3810_0 = v_3811_0 | v_10164_0;
  assign v_3811_0 = v_589_0 ? v_3812_0 : 3'h0;
  assign v_3813_0 = v_3814_0 | v_3815_0;
  assign v_3814_0 = v_589_0 | v_601_0;
  assign v_3815_0 = v_607_0 | v_26_0;
  assign v_3816_0 = v_3817_0 | v_10161_0;
  assign v_3817_0 = v_3818_0 | v_10160_0;
  assign v_3818_0 = v_589_0 ? v_3819_0 : 3'h0;
  assign v_3820_0 = v_3821_0 | v_3822_0;
  assign v_3821_0 = v_589_0 | v_601_0;
  assign v_3822_0 = v_607_0 | v_26_0;
  assign v_3823_0 = v_3824_0 | v_10157_0;
  assign v_3824_0 = v_3825_0 | v_10156_0;
  assign v_3825_0 = v_589_0 ? v_3826_0 : 3'h0;
  assign v_3827_0 = v_3828_0 | v_3829_0;
  assign v_3828_0 = v_589_0 | v_601_0;
  assign v_3829_0 = v_607_0 | v_26_0;
  assign v_3830_0 = v_3831_0 | v_10153_0;
  assign v_3831_0 = v_3832_0 | v_10152_0;
  assign v_3832_0 = v_589_0 ? v_3833_0 : 3'h0;
  assign v_3834_0 = v_3835_0 | v_3836_0;
  assign v_3835_0 = v_589_0 | v_601_0;
  assign v_3836_0 = v_607_0 | v_26_0;
  assign v_3837_0 = v_3838_0 | v_10149_0;
  assign v_3838_0 = v_3839_0 | v_10148_0;
  assign v_3839_0 = v_589_0 ? v_3840_0 : 3'h0;
  assign v_3841_0 = v_3842_0 | v_3843_0;
  assign v_3842_0 = v_589_0 | v_601_0;
  assign v_3843_0 = v_607_0 | v_26_0;
  assign v_3844_0 = v_3845_0 | v_10145_0;
  assign v_3845_0 = v_3846_0 | v_10144_0;
  assign v_3846_0 = v_589_0 ? v_3847_0 : 3'h0;
  assign v_3848_0 = v_3849_0 | v_3850_0;
  assign v_3849_0 = v_589_0 | v_601_0;
  assign v_3850_0 = v_607_0 | v_26_0;
  assign v_3851_0 = v_3852_0 | v_10141_0;
  assign v_3852_0 = v_3853_0 | v_10140_0;
  assign v_3853_0 = v_589_0 ? v_3854_0 : 3'h0;
  assign v_3855_0 = v_3856_0 | v_3857_0;
  assign v_3856_0 = v_589_0 | v_601_0;
  assign v_3857_0 = v_607_0 | v_26_0;
  assign v_3858_0 = v_3859_0 | v_10137_0;
  assign v_3859_0 = v_3860_0 | v_10136_0;
  assign v_3860_0 = v_589_0 ? v_3861_0 : 3'h0;
  assign v_3862_0 = v_3863_0 | v_3864_0;
  assign v_3863_0 = v_589_0 | v_601_0;
  assign v_3864_0 = v_607_0 | v_26_0;
  assign v_3865_0 = v_3866_0 | v_10133_0;
  assign v_3866_0 = v_3867_0 | v_10132_0;
  assign v_3867_0 = v_589_0 ? v_3868_0 : 3'h0;
  assign v_3869_0 = v_3870_0 | v_3871_0;
  assign v_3870_0 = v_589_0 | v_601_0;
  assign v_3871_0 = v_607_0 | v_26_0;
  assign v_3872_0 = v_3873_0 | v_10129_0;
  assign v_3873_0 = v_3874_0 | v_10128_0;
  assign v_3874_0 = v_589_0 ? v_3875_0 : 3'h0;
  assign v_3876_0 = v_3877_0 | v_3878_0;
  assign v_3877_0 = v_589_0 | v_601_0;
  assign v_3878_0 = v_607_0 | v_26_0;
  assign v_3879_0 = v_3880_0 | v_10125_0;
  assign v_3880_0 = v_3881_0 | v_10124_0;
  assign v_3881_0 = v_589_0 ? v_3882_0 : 3'h0;
  assign v_3883_0 = v_3884_0 | v_3885_0;
  assign v_3884_0 = v_589_0 | v_601_0;
  assign v_3885_0 = v_607_0 | v_26_0;
  assign v_3886_0 = v_3887_0 | v_10121_0;
  assign v_3887_0 = v_3888_0 | v_10120_0;
  assign v_3888_0 = v_589_0 ? v_3889_0 : 3'h0;
  assign v_3890_0 = v_3891_0 | v_3892_0;
  assign v_3891_0 = v_589_0 | v_601_0;
  assign v_3892_0 = v_607_0 | v_26_0;
  assign v_3893_0 = v_3894_0 | v_10117_0;
  assign v_3894_0 = v_3895_0 | v_10116_0;
  assign v_3895_0 = v_589_0 ? v_3896_0 : 3'h0;
  assign v_3897_0 = v_3898_0 | v_3899_0;
  assign v_3898_0 = v_589_0 | v_601_0;
  assign v_3899_0 = v_607_0 | v_26_0;
  assign v_3900_0 = v_3901_0 | v_10113_0;
  assign v_3901_0 = v_3902_0 | v_10112_0;
  assign v_3902_0 = v_589_0 ? v_3903_0 : 3'h0;
  assign v_3904_0 = v_3905_0 | v_3906_0;
  assign v_3905_0 = v_589_0 | v_601_0;
  assign v_3906_0 = v_607_0 | v_26_0;
  assign v_3907_0 = v_3908_0 | v_10109_0;
  assign v_3908_0 = v_3909_0 | v_10108_0;
  assign v_3909_0 = v_589_0 ? v_3910_0 : 3'h0;
  assign v_3911_0 = v_3912_0 | v_3913_0;
  assign v_3912_0 = v_589_0 | v_601_0;
  assign v_3913_0 = v_607_0 | v_26_0;
  assign v_3914_0 = v_3915_0 | v_10105_0;
  assign v_3915_0 = v_3916_0 | v_10104_0;
  assign v_3916_0 = v_589_0 ? v_3917_0 : 3'h0;
  assign v_3918_0 = v_3919_0 | v_3920_0;
  assign v_3919_0 = v_589_0 | v_601_0;
  assign v_3920_0 = v_607_0 | v_26_0;
  assign v_3921_0 = v_3922_0 | v_10101_0;
  assign v_3922_0 = v_3923_0 | v_10100_0;
  assign v_3923_0 = v_589_0 ? v_3924_0 : 3'h0;
  assign v_3925_0 = v_3926_0 | v_3927_0;
  assign v_3926_0 = v_589_0 | v_601_0;
  assign v_3927_0 = v_607_0 | v_26_0;
  assign v_3928_0 = v_3929_0 | v_10097_0;
  assign v_3929_0 = v_3930_0 | v_10096_0;
  assign v_3930_0 = v_589_0 ? v_3931_0 : 3'h0;
  assign v_3932_0 = v_3933_0 | v_3934_0;
  assign v_3933_0 = v_589_0 | v_601_0;
  assign v_3934_0 = v_607_0 | v_26_0;
  assign v_3935_0 = v_3936_0 | v_10093_0;
  assign v_3936_0 = v_3937_0 | v_10092_0;
  assign v_3937_0 = v_589_0 ? v_3938_0 : 3'h0;
  assign v_3939_0 = v_3940_0 | v_3941_0;
  assign v_3940_0 = v_589_0 | v_601_0;
  assign v_3941_0 = v_607_0 | v_26_0;
  assign v_3942_0 = v_3943_0 | v_10089_0;
  assign v_3943_0 = v_3944_0 | v_10088_0;
  assign v_3944_0 = v_589_0 ? v_3945_0 : 3'h0;
  assign v_3946_0 = v_3947_0 | v_3948_0;
  assign v_3947_0 = v_589_0 | v_601_0;
  assign v_3948_0 = v_607_0 | v_26_0;
  assign v_3949_0 = v_3950_0 | v_10085_0;
  assign v_3950_0 = v_3951_0 | v_10084_0;
  assign v_3951_0 = v_589_0 ? v_3952_0 : 3'h0;
  assign v_3953_0 = v_3954_0 | v_3955_0;
  assign v_3954_0 = v_589_0 | v_601_0;
  assign v_3955_0 = v_607_0 | v_26_0;
  assign v_3956_0 = v_3957_0 | v_10081_0;
  assign v_3957_0 = v_3958_0 | v_10080_0;
  assign v_3958_0 = v_589_0 ? v_3959_0 : 3'h0;
  assign v_3960_0 = v_3961_0 | v_3962_0;
  assign v_3961_0 = v_589_0 | v_601_0;
  assign v_3962_0 = v_607_0 | v_26_0;
  assign v_3963_0 = v_3964_0 | v_10077_0;
  assign v_3964_0 = v_3965_0 | v_10076_0;
  assign v_3965_0 = v_589_0 ? v_3966_0 : 3'h0;
  assign v_3967_0 = v_3968_0 | v_3969_0;
  assign v_3968_0 = v_589_0 | v_601_0;
  assign v_3969_0 = v_607_0 | v_26_0;
  assign v_3970_0 = v_3971_0 | v_10073_0;
  assign v_3971_0 = v_3972_0 | v_10072_0;
  assign v_3972_0 = v_589_0 ? v_3973_0 : 3'h0;
  assign v_3974_0 = v_3975_0 | v_3976_0;
  assign v_3975_0 = v_589_0 | v_601_0;
  assign v_3976_0 = v_607_0 | v_26_0;
  assign v_3977_0 = v_3978_0 | v_10069_0;
  assign v_3978_0 = v_3979_0 | v_10068_0;
  assign v_3979_0 = v_589_0 ? v_3980_0 : 3'h0;
  assign v_3981_0 = v_3982_0 | v_3983_0;
  assign v_3982_0 = v_589_0 | v_601_0;
  assign v_3983_0 = v_607_0 | v_26_0;
  assign v_3984_0 = v_3985_0 | v_10065_0;
  assign v_3985_0 = v_3986_0 | v_10064_0;
  assign v_3986_0 = v_589_0 ? v_3987_0 : 3'h0;
  assign v_3988_0 = v_3989_0 | v_3990_0;
  assign v_3989_0 = v_589_0 | v_601_0;
  assign v_3990_0 = v_607_0 | v_26_0;
  assign v_3991_0 = v_3992_0 | v_10061_0;
  assign v_3992_0 = v_3993_0 | v_10060_0;
  assign v_3993_0 = v_589_0 ? v_3994_0 : 3'h0;
  assign v_3995_0 = v_3996_0 | v_3997_0;
  assign v_3996_0 = v_589_0 | v_601_0;
  assign v_3997_0 = v_607_0 | v_26_0;
  assign v_3998_0 = v_3999_0 | v_10057_0;
  assign v_3999_0 = v_4000_0 | v_10056_0;
  assign v_4000_0 = v_589_0 ? v_4001_0 : 3'h0;
  assign v_4002_0 = v_4003_0 | v_4004_0;
  assign v_4003_0 = v_589_0 | v_601_0;
  assign v_4004_0 = v_607_0 | v_26_0;
  assign v_4005_0 = v_4006_0 | v_10053_0;
  assign v_4006_0 = v_4007_0 | v_10052_0;
  assign v_4007_0 = v_589_0 ? v_4008_0 : 3'h0;
  assign v_4009_0 = v_4010_0 | v_4011_0;
  assign v_4010_0 = v_589_0 | v_601_0;
  assign v_4011_0 = v_607_0 | v_26_0;
  assign v_4012_0 = v_4013_0 | v_10049_0;
  assign v_4013_0 = v_4014_0 | v_10048_0;
  assign v_4014_0 = v_589_0 ? v_4015_0 : 3'h0;
  assign v_4016_0 = v_4017_0 | v_4018_0;
  assign v_4017_0 = v_589_0 | v_601_0;
  assign v_4018_0 = v_607_0 | v_26_0;
  assign v_4019_0 = v_4020_0 | v_10045_0;
  assign v_4020_0 = v_4021_0 | v_10044_0;
  assign v_4021_0 = v_589_0 ? v_4022_0 : 3'h0;
  assign v_4023_0 = v_4024_0 | v_4025_0;
  assign v_4024_0 = v_589_0 | v_601_0;
  assign v_4025_0 = v_607_0 | v_26_0;
  assign v_4026_0 = v_4027_0 | v_10041_0;
  assign v_4027_0 = v_4028_0 | v_10040_0;
  assign v_4028_0 = v_589_0 ? v_4029_0 : 3'h0;
  assign v_4030_0 = v_4031_0 | v_4032_0;
  assign v_4031_0 = v_589_0 | v_601_0;
  assign v_4032_0 = v_607_0 | v_26_0;
  assign v_4033_0 = v_4034_0 | v_10037_0;
  assign v_4034_0 = v_4035_0 | v_10036_0;
  assign v_4035_0 = v_589_0 ? v_4036_0 : 3'h0;
  assign v_4037_0 = v_4038_0 | v_4039_0;
  assign v_4038_0 = v_589_0 | v_601_0;
  assign v_4039_0 = v_607_0 | v_26_0;
  assign v_4040_0 = v_4041_0 | v_10033_0;
  assign v_4041_0 = v_4042_0 | v_10032_0;
  assign v_4042_0 = v_589_0 ? v_4043_0 : 3'h0;
  assign v_4044_0 = v_4045_0 | v_4046_0;
  assign v_4045_0 = v_589_0 | v_601_0;
  assign v_4046_0 = v_607_0 | v_26_0;
  assign v_4047_0 = v_4048_0 | v_10029_0;
  assign v_4048_0 = v_4049_0 | v_10028_0;
  assign v_4049_0 = v_589_0 ? v_4050_0 : 3'h0;
  assign v_4051_0 = v_4052_0 | v_4053_0;
  assign v_4052_0 = v_589_0 | v_601_0;
  assign v_4053_0 = v_607_0 | v_26_0;
  assign v_4054_0 = v_4055_0 | v_10025_0;
  assign v_4055_0 = v_4056_0 | v_10024_0;
  assign v_4056_0 = v_589_0 ? v_4057_0 : 3'h0;
  assign v_4058_0 = v_4059_0 | v_4060_0;
  assign v_4059_0 = v_589_0 | v_601_0;
  assign v_4060_0 = v_607_0 | v_26_0;
  assign v_4061_0 = v_4062_0 | v_10021_0;
  assign v_4062_0 = v_4063_0 | v_10020_0;
  assign v_4063_0 = v_589_0 ? v_4064_0 : 3'h0;
  assign v_4065_0 = v_4066_0 | v_4067_0;
  assign v_4066_0 = v_589_0 | v_601_0;
  assign v_4067_0 = v_607_0 | v_26_0;
  assign v_4068_0 = v_4069_0 | v_10017_0;
  assign v_4069_0 = v_4070_0 | v_10016_0;
  assign v_4070_0 = v_589_0 ? v_4071_0 : 3'h0;
  assign v_4072_0 = v_4073_0 | v_4074_0;
  assign v_4073_0 = v_589_0 | v_601_0;
  assign v_4074_0 = v_607_0 | v_26_0;
  assign v_4075_0 = v_4076_0 | v_10013_0;
  assign v_4076_0 = v_4077_0 | v_10012_0;
  assign v_4077_0 = v_589_0 ? v_4078_0 : 3'h0;
  assign v_4079_0 = v_4080_0 | v_4081_0;
  assign v_4080_0 = v_589_0 | v_601_0;
  assign v_4081_0 = v_607_0 | v_26_0;
  assign v_4082_0 = v_4083_0 | v_10009_0;
  assign v_4083_0 = v_4084_0 | v_10008_0;
  assign v_4084_0 = v_589_0 ? v_4085_0 : 3'h0;
  assign v_4086_0 = v_4087_0 | v_4088_0;
  assign v_4087_0 = v_589_0 | v_601_0;
  assign v_4088_0 = v_607_0 | v_26_0;
  assign v_4089_0 = v_4090_0 | v_10005_0;
  assign v_4090_0 = v_4091_0 | v_10004_0;
  assign v_4091_0 = v_589_0 ? v_4092_0 : 3'h0;
  assign v_4093_0 = v_4094_0 | v_4095_0;
  assign v_4094_0 = v_589_0 | v_601_0;
  assign v_4095_0 = v_607_0 | v_26_0;
  assign v_4096_0 = v_4097_0 | v_10001_0;
  assign v_4097_0 = v_4098_0 | v_10000_0;
  assign v_4098_0 = v_589_0 ? v_4099_0 : 3'h0;
  assign v_4100_0 = v_4101_0 | v_4102_0;
  assign v_4101_0 = v_589_0 | v_601_0;
  assign v_4102_0 = v_607_0 | v_26_0;
  assign v_4103_0 = v_4104_0 | v_9997_0;
  assign v_4104_0 = v_4105_0 | v_9996_0;
  assign v_4105_0 = v_589_0 ? v_4106_0 : 3'h0;
  assign v_4107_0 = v_4108_0 | v_4109_0;
  assign v_4108_0 = v_589_0 | v_601_0;
  assign v_4109_0 = v_607_0 | v_26_0;
  assign v_4110_0 = v_4111_0 | v_9993_0;
  assign v_4111_0 = v_4112_0 | v_9992_0;
  assign v_4112_0 = v_589_0 ? v_4113_0 : 3'h0;
  assign v_4114_0 = v_4115_0 | v_4116_0;
  assign v_4115_0 = v_589_0 | v_601_0;
  assign v_4116_0 = v_607_0 | v_26_0;
  assign v_4117_0 = v_4118_0 | v_9989_0;
  assign v_4118_0 = v_4119_0 | v_9988_0;
  assign v_4119_0 = v_589_0 ? v_4120_0 : 3'h0;
  assign v_4121_0 = v_4122_0 | v_4123_0;
  assign v_4122_0 = v_589_0 | v_601_0;
  assign v_4123_0 = v_607_0 | v_26_0;
  assign v_4124_0 = v_4125_0 | v_9985_0;
  assign v_4125_0 = v_4126_0 | v_9984_0;
  assign v_4126_0 = v_589_0 ? v_4127_0 : 3'h0;
  assign v_4128_0 = v_4129_0 | v_4130_0;
  assign v_4129_0 = v_589_0 | v_601_0;
  assign v_4130_0 = v_607_0 | v_26_0;
  assign v_4131_0 = v_4132_0 | v_9981_0;
  assign v_4132_0 = v_4133_0 | v_9980_0;
  assign v_4133_0 = v_589_0 ? v_4134_0 : 3'h0;
  assign v_4135_0 = v_4136_0 | v_4137_0;
  assign v_4136_0 = v_589_0 | v_601_0;
  assign v_4137_0 = v_607_0 | v_26_0;
  assign v_4138_0 = v_4139_0 | v_9977_0;
  assign v_4139_0 = v_4140_0 | v_9976_0;
  assign v_4140_0 = v_589_0 ? v_4141_0 : 3'h0;
  assign v_4142_0 = v_4143_0 | v_4144_0;
  assign v_4143_0 = v_589_0 | v_601_0;
  assign v_4144_0 = v_607_0 | v_26_0;
  assign v_4145_0 = v_4146_0 | v_9973_0;
  assign v_4146_0 = v_4147_0 | v_9972_0;
  assign v_4147_0 = v_589_0 ? v_4148_0 : 3'h0;
  assign v_4149_0 = v_4150_0 | v_4151_0;
  assign v_4150_0 = v_589_0 | v_601_0;
  assign v_4151_0 = v_607_0 | v_26_0;
  assign v_4152_0 = v_4153_0 | v_9969_0;
  assign v_4153_0 = v_4154_0 | v_9968_0;
  assign v_4154_0 = v_589_0 ? v_4155_0 : 3'h0;
  assign v_4156_0 = v_4157_0 | v_4158_0;
  assign v_4157_0 = v_589_0 | v_601_0;
  assign v_4158_0 = v_607_0 | v_26_0;
  assign v_4159_0 = v_4160_0 | v_9965_0;
  assign v_4160_0 = v_4161_0 | v_9964_0;
  assign v_4161_0 = v_589_0 ? v_4162_0 : 3'h0;
  assign v_4163_0 = v_4164_0 | v_4165_0;
  assign v_4164_0 = v_589_0 | v_601_0;
  assign v_4165_0 = v_607_0 | v_26_0;
  assign v_4166_0 = v_4167_0 | v_9961_0;
  assign v_4167_0 = v_4168_0 | v_9960_0;
  assign v_4168_0 = v_589_0 ? v_4169_0 : 3'h0;
  assign v_4170_0 = v_4171_0 | v_4172_0;
  assign v_4171_0 = v_589_0 | v_601_0;
  assign v_4172_0 = v_607_0 | v_26_0;
  assign v_4173_0 = v_4174_0 | v_9957_0;
  assign v_4174_0 = v_4175_0 | v_9956_0;
  assign v_4175_0 = v_589_0 ? v_4176_0 : 3'h0;
  assign v_4177_0 = v_4178_0 | v_4179_0;
  assign v_4178_0 = v_589_0 | v_601_0;
  assign v_4179_0 = v_607_0 | v_26_0;
  assign v_4180_0 = v_4181_0 | v_9953_0;
  assign v_4181_0 = v_4182_0 | v_9952_0;
  assign v_4182_0 = v_589_0 ? v_4183_0 : 3'h0;
  assign v_4184_0 = v_4185_0 | v_4186_0;
  assign v_4185_0 = v_589_0 | v_601_0;
  assign v_4186_0 = v_607_0 | v_26_0;
  assign v_4187_0 = v_4188_0 | v_9949_0;
  assign v_4188_0 = v_4189_0 | v_9948_0;
  assign v_4189_0 = v_589_0 ? v_4190_0 : 3'h0;
  assign v_4191_0 = v_4192_0 | v_4193_0;
  assign v_4192_0 = v_589_0 | v_601_0;
  assign v_4193_0 = v_607_0 | v_26_0;
  assign v_4194_0 = v_4195_0 | v_9945_0;
  assign v_4195_0 = v_4196_0 | v_9944_0;
  assign v_4196_0 = v_589_0 ? v_4197_0 : 3'h0;
  assign v_4198_0 = v_4199_0 | v_4200_0;
  assign v_4199_0 = v_589_0 | v_601_0;
  assign v_4200_0 = v_607_0 | v_26_0;
  assign v_4201_0 = v_4202_0 | v_9941_0;
  assign v_4202_0 = v_4203_0 | v_9940_0;
  assign v_4203_0 = v_589_0 ? v_4204_0 : 3'h0;
  assign v_4205_0 = v_4206_0 | v_4207_0;
  assign v_4206_0 = v_589_0 | v_601_0;
  assign v_4207_0 = v_607_0 | v_26_0;
  assign v_4208_0 = v_4209_0 | v_9937_0;
  assign v_4209_0 = v_4210_0 | v_9936_0;
  assign v_4210_0 = v_589_0 ? v_4211_0 : 3'h0;
  assign v_4212_0 = v_4213_0 | v_4214_0;
  assign v_4213_0 = v_589_0 | v_601_0;
  assign v_4214_0 = v_607_0 | v_26_0;
  assign v_4215_0 = v_4216_0 | v_9933_0;
  assign v_4216_0 = v_4217_0 | v_9932_0;
  assign v_4217_0 = v_589_0 ? v_4218_0 : 3'h0;
  assign v_4219_0 = v_4220_0 | v_4221_0;
  assign v_4220_0 = v_589_0 | v_601_0;
  assign v_4221_0 = v_607_0 | v_26_0;
  assign v_4222_0 = v_4223_0 | v_9929_0;
  assign v_4223_0 = v_4224_0 | v_9928_0;
  assign v_4224_0 = v_589_0 ? v_4225_0 : 3'h0;
  assign v_4226_0 = v_4227_0 | v_4228_0;
  assign v_4227_0 = v_589_0 | v_601_0;
  assign v_4228_0 = v_607_0 | v_26_0;
  assign v_4229_0 = v_4230_0 | v_9925_0;
  assign v_4230_0 = v_4231_0 | v_9924_0;
  assign v_4231_0 = v_589_0 ? v_4232_0 : 3'h0;
  assign v_4233_0 = v_4234_0 | v_4235_0;
  assign v_4234_0 = v_589_0 | v_601_0;
  assign v_4235_0 = v_607_0 | v_26_0;
  assign v_4236_0 = v_4237_0 | v_9921_0;
  assign v_4237_0 = v_4238_0 | v_9920_0;
  assign v_4238_0 = v_589_0 ? v_4239_0 : 3'h0;
  assign v_4240_0 = v_4241_0 | v_4242_0;
  assign v_4241_0 = v_589_0 | v_601_0;
  assign v_4242_0 = v_607_0 | v_26_0;
  assign v_4243_0 = v_4244_0 | v_9917_0;
  assign v_4244_0 = v_4245_0 | v_9916_0;
  assign v_4245_0 = v_589_0 ? v_4246_0 : 3'h0;
  assign v_4247_0 = v_4248_0 | v_4249_0;
  assign v_4248_0 = v_589_0 | v_601_0;
  assign v_4249_0 = v_607_0 | v_26_0;
  assign v_4250_0 = v_4251_0 | v_9913_0;
  assign v_4251_0 = v_4252_0 | v_9912_0;
  assign v_4252_0 = v_589_0 ? v_4253_0 : 3'h0;
  assign v_4254_0 = v_4255_0 | v_4256_0;
  assign v_4255_0 = v_589_0 | v_601_0;
  assign v_4256_0 = v_607_0 | v_26_0;
  assign v_4257_0 = v_4258_0 | v_9909_0;
  assign v_4258_0 = v_4259_0 | v_9908_0;
  assign v_4259_0 = v_589_0 ? v_4260_0 : 3'h0;
  assign v_4261_0 = v_4262_0 | v_4263_0;
  assign v_4262_0 = v_589_0 | v_601_0;
  assign v_4263_0 = v_607_0 | v_26_0;
  assign v_4264_0 = v_4265_0 | v_9905_0;
  assign v_4265_0 = v_4266_0 | v_9904_0;
  assign v_4266_0 = v_589_0 ? v_4267_0 : 3'h0;
  assign v_4268_0 = v_4269_0 | v_4270_0;
  assign v_4269_0 = v_589_0 | v_601_0;
  assign v_4270_0 = v_607_0 | v_26_0;
  assign v_4271_0 = v_4272_0 | v_9901_0;
  assign v_4272_0 = v_4273_0 | v_9900_0;
  assign v_4273_0 = v_589_0 ? v_4274_0 : 3'h0;
  assign v_4275_0 = v_4276_0 | v_4277_0;
  assign v_4276_0 = v_589_0 | v_601_0;
  assign v_4277_0 = v_607_0 | v_26_0;
  assign v_4278_0 = v_4279_0 | v_9897_0;
  assign v_4279_0 = v_4280_0 | v_9896_0;
  assign v_4280_0 = v_589_0 ? v_4281_0 : 3'h0;
  assign v_4282_0 = v_4283_0 | v_4284_0;
  assign v_4283_0 = v_589_0 | v_601_0;
  assign v_4284_0 = v_607_0 | v_26_0;
  assign v_4285_0 = v_4286_0 | v_9893_0;
  assign v_4286_0 = v_4287_0 | v_9892_0;
  assign v_4287_0 = v_589_0 ? v_4288_0 : 3'h0;
  assign v_4289_0 = v_4290_0 | v_4291_0;
  assign v_4290_0 = v_589_0 | v_601_0;
  assign v_4291_0 = v_607_0 | v_26_0;
  assign v_4292_0 = v_4293_0 | v_9889_0;
  assign v_4293_0 = v_4294_0 | v_9888_0;
  assign v_4294_0 = v_589_0 ? v_4295_0 : 3'h0;
  assign v_4296_0 = v_4297_0 | v_4298_0;
  assign v_4297_0 = v_589_0 | v_601_0;
  assign v_4298_0 = v_607_0 | v_26_0;
  assign v_4299_0 = v_4300_0 | v_9885_0;
  assign v_4300_0 = v_4301_0 | v_9884_0;
  assign v_4301_0 = v_589_0 ? v_4302_0 : 3'h0;
  assign v_4303_0 = v_4304_0 | v_4305_0;
  assign v_4304_0 = v_589_0 | v_601_0;
  assign v_4305_0 = v_607_0 | v_26_0;
  assign v_4306_0 = v_4307_0 | v_9881_0;
  assign v_4307_0 = v_4308_0 | v_9880_0;
  assign v_4308_0 = v_589_0 ? v_4309_0 : 3'h0;
  assign v_4310_0 = v_4311_0 | v_4312_0;
  assign v_4311_0 = v_589_0 | v_601_0;
  assign v_4312_0 = v_607_0 | v_26_0;
  assign v_4313_0 = v_4314_0 | v_9877_0;
  assign v_4314_0 = v_4315_0 | v_9876_0;
  assign v_4315_0 = v_589_0 ? v_4316_0 : 3'h0;
  assign v_4317_0 = v_4318_0 | v_4319_0;
  assign v_4318_0 = v_589_0 | v_601_0;
  assign v_4319_0 = v_607_0 | v_26_0;
  assign v_4320_0 = v_4321_0 | v_9873_0;
  assign v_4321_0 = v_4322_0 | v_9872_0;
  assign v_4322_0 = v_589_0 ? v_4323_0 : 3'h0;
  assign v_4324_0 = v_4325_0 | v_4326_0;
  assign v_4325_0 = v_589_0 | v_601_0;
  assign v_4326_0 = v_607_0 | v_26_0;
  assign v_4327_0 = v_4328_0 | v_9869_0;
  assign v_4328_0 = v_4329_0 | v_9868_0;
  assign v_4329_0 = v_589_0 ? v_4330_0 : 3'h0;
  assign v_4331_0 = v_4332_0 | v_4333_0;
  assign v_4332_0 = v_589_0 | v_601_0;
  assign v_4333_0 = v_607_0 | v_26_0;
  assign v_4334_0 = v_4335_0 | v_9865_0;
  assign v_4335_0 = v_4336_0 | v_9864_0;
  assign v_4336_0 = v_589_0 ? v_4337_0 : 3'h0;
  assign v_4338_0 = v_4339_0 | v_4340_0;
  assign v_4339_0 = v_589_0 | v_601_0;
  assign v_4340_0 = v_607_0 | v_26_0;
  assign v_4341_0 = v_4342_0 | v_9861_0;
  assign v_4342_0 = v_4343_0 | v_9860_0;
  assign v_4343_0 = v_589_0 ? v_4344_0 : 3'h0;
  assign v_4345_0 = v_4346_0 | v_4347_0;
  assign v_4346_0 = v_589_0 | v_601_0;
  assign v_4347_0 = v_607_0 | v_26_0;
  assign v_4348_0 = v_4349_0 | v_9857_0;
  assign v_4349_0 = v_4350_0 | v_9856_0;
  assign v_4350_0 = v_589_0 ? v_4351_0 : 3'h0;
  assign v_4352_0 = v_4353_0 | v_4354_0;
  assign v_4353_0 = v_589_0 | v_601_0;
  assign v_4354_0 = v_607_0 | v_26_0;
  assign v_4355_0 = v_4356_0 | v_9853_0;
  assign v_4356_0 = v_4357_0 | v_9852_0;
  assign v_4357_0 = v_589_0 ? v_4358_0 : 3'h0;
  assign v_4359_0 = v_4360_0 | v_4361_0;
  assign v_4360_0 = v_589_0 | v_601_0;
  assign v_4361_0 = v_607_0 | v_26_0;
  assign v_4362_0 = v_4363_0 | v_9849_0;
  assign v_4363_0 = v_4364_0 | v_9848_0;
  assign v_4364_0 = v_589_0 ? v_4365_0 : 3'h0;
  assign v_4366_0 = v_4367_0 | v_4368_0;
  assign v_4367_0 = v_589_0 | v_601_0;
  assign v_4368_0 = v_607_0 | v_26_0;
  assign v_4369_0 = v_4370_0 | v_9845_0;
  assign v_4370_0 = v_4371_0 | v_9844_0;
  assign v_4371_0 = v_589_0 ? v_4372_0 : 3'h0;
  assign v_4373_0 = v_4374_0 | v_4375_0;
  assign v_4374_0 = v_589_0 | v_601_0;
  assign v_4375_0 = v_607_0 | v_26_0;
  assign v_4376_0 = v_4377_0 | v_9841_0;
  assign v_4377_0 = v_4378_0 | v_9840_0;
  assign v_4378_0 = v_589_0 ? v_4379_0 : 3'h0;
  assign v_4380_0 = v_4381_0 | v_4382_0;
  assign v_4381_0 = v_589_0 | v_601_0;
  assign v_4382_0 = v_607_0 | v_26_0;
  assign v_4383_0 = v_4384_0 | v_9837_0;
  assign v_4384_0 = v_4385_0 | v_9836_0;
  assign v_4385_0 = v_589_0 ? v_4386_0 : 3'h0;
  assign v_4387_0 = v_4388_0 | v_4389_0;
  assign v_4388_0 = v_589_0 | v_601_0;
  assign v_4389_0 = v_607_0 | v_26_0;
  assign v_4390_0 = v_4391_0 | v_9833_0;
  assign v_4391_0 = v_4392_0 | v_9832_0;
  assign v_4392_0 = v_589_0 ? v_4393_0 : 3'h0;
  assign v_4394_0 = v_4395_0 | v_4396_0;
  assign v_4395_0 = v_589_0 | v_601_0;
  assign v_4396_0 = v_607_0 | v_26_0;
  assign v_4397_0 = v_4398_0 | v_9829_0;
  assign v_4398_0 = v_4399_0 | v_9828_0;
  assign v_4399_0 = v_589_0 ? v_4400_0 : 3'h0;
  assign v_4401_0 = v_4402_0 | v_4403_0;
  assign v_4402_0 = v_589_0 | v_601_0;
  assign v_4403_0 = v_607_0 | v_26_0;
  assign v_4404_0 = v_4405_0 | v_9825_0;
  assign v_4405_0 = v_4406_0 | v_9824_0;
  assign v_4406_0 = v_589_0 ? v_4407_0 : 3'h0;
  assign v_4408_0 = v_4409_0 | v_4410_0;
  assign v_4409_0 = v_589_0 | v_601_0;
  assign v_4410_0 = v_607_0 | v_26_0;
  assign v_4411_0 = v_4412_0 | v_9821_0;
  assign v_4412_0 = v_4413_0 | v_9820_0;
  assign v_4413_0 = v_589_0 ? v_4414_0 : 3'h0;
  assign v_4415_0 = v_4416_0 | v_4417_0;
  assign v_4416_0 = v_589_0 | v_601_0;
  assign v_4417_0 = v_607_0 | v_26_0;
  assign v_4418_0 = v_4419_0 | v_9817_0;
  assign v_4419_0 = v_4420_0 | v_9816_0;
  assign v_4420_0 = v_589_0 ? v_4421_0 : 3'h0;
  assign v_4422_0 = v_4423_0 | v_4424_0;
  assign v_4423_0 = v_589_0 | v_601_0;
  assign v_4424_0 = v_607_0 | v_26_0;
  assign v_4425_0 = v_4426_0 | v_9813_0;
  assign v_4426_0 = v_4427_0 | v_9812_0;
  assign v_4427_0 = v_589_0 ? v_4428_0 : 3'h0;
  assign v_4429_0 = v_4430_0 | v_4431_0;
  assign v_4430_0 = v_589_0 | v_601_0;
  assign v_4431_0 = v_607_0 | v_26_0;
  assign v_4432_0 = v_4433_0 | v_9809_0;
  assign v_4433_0 = v_4434_0 | v_9808_0;
  assign v_4434_0 = v_589_0 ? v_4435_0 : 3'h0;
  assign v_4436_0 = v_4437_0 | v_4438_0;
  assign v_4437_0 = v_589_0 | v_601_0;
  assign v_4438_0 = v_607_0 | v_26_0;
  assign v_4439_0 = v_4440_0 | v_9805_0;
  assign v_4440_0 = v_4441_0 | v_9804_0;
  assign v_4441_0 = v_589_0 ? v_4442_0 : 3'h0;
  assign v_4443_0 = v_4444_0 | v_4445_0;
  assign v_4444_0 = v_589_0 | v_601_0;
  assign v_4445_0 = v_607_0 | v_26_0;
  assign v_4446_0 = v_4447_0 | v_9801_0;
  assign v_4447_0 = v_4448_0 | v_9800_0;
  assign v_4448_0 = v_589_0 ? v_4449_0 : 3'h0;
  assign v_4450_0 = v_4451_0 | v_4452_0;
  assign v_4451_0 = v_589_0 | v_601_0;
  assign v_4452_0 = v_607_0 | v_26_0;
  assign v_4453_0 = v_4454_0 | v_9797_0;
  assign v_4454_0 = v_4455_0 | v_9796_0;
  assign v_4455_0 = v_589_0 ? v_4456_0 : 3'h0;
  assign v_4457_0 = v_4458_0 | v_4459_0;
  assign v_4458_0 = v_589_0 | v_601_0;
  assign v_4459_0 = v_607_0 | v_26_0;
  assign v_4460_0 = v_4461_0 | v_9793_0;
  assign v_4461_0 = v_4462_0 | v_9792_0;
  assign v_4462_0 = v_589_0 ? v_4463_0 : 3'h0;
  assign v_4464_0 = v_4465_0 | v_4466_0;
  assign v_4465_0 = v_589_0 | v_601_0;
  assign v_4466_0 = v_607_0 | v_26_0;
  assign v_4467_0 = v_4468_0 | v_9789_0;
  assign v_4468_0 = v_4469_0 | v_9788_0;
  assign v_4469_0 = v_589_0 ? v_4470_0 : 3'h0;
  assign v_4471_0 = v_4472_0 | v_4473_0;
  assign v_4472_0 = v_589_0 | v_601_0;
  assign v_4473_0 = v_607_0 | v_26_0;
  assign v_4474_0 = v_4475_0 | v_9785_0;
  assign v_4475_0 = v_4476_0 | v_9784_0;
  assign v_4476_0 = v_589_0 ? v_4477_0 : 3'h0;
  assign v_4478_0 = v_4479_0 | v_4480_0;
  assign v_4479_0 = v_589_0 | v_601_0;
  assign v_4480_0 = v_607_0 | v_26_0;
  assign v_4481_0 = v_4482_0 | v_9781_0;
  assign v_4482_0 = v_4483_0 | v_9780_0;
  assign v_4483_0 = v_589_0 ? v_4484_0 : 3'h0;
  assign v_4485_0 = v_4486_0 | v_4487_0;
  assign v_4486_0 = v_589_0 | v_601_0;
  assign v_4487_0 = v_607_0 | v_26_0;
  assign v_4488_0 = v_4489_0 | v_9777_0;
  assign v_4489_0 = v_4490_0 | v_9776_0;
  assign v_4490_0 = v_589_0 ? v_4491_0 : 3'h0;
  assign v_4492_0 = v_4493_0 | v_4494_0;
  assign v_4493_0 = v_589_0 | v_601_0;
  assign v_4494_0 = v_607_0 | v_26_0;
  assign v_4495_0 = v_4496_0 | v_9773_0;
  assign v_4496_0 = v_4497_0 | v_9772_0;
  assign v_4497_0 = v_589_0 ? v_4498_0 : 3'h0;
  assign v_4499_0 = v_4500_0 | v_4501_0;
  assign v_4500_0 = v_589_0 | v_601_0;
  assign v_4501_0 = v_607_0 | v_26_0;
  assign v_4502_0 = v_4503_0 | v_9769_0;
  assign v_4503_0 = v_4504_0 | v_9768_0;
  assign v_4504_0 = v_589_0 ? v_4505_0 : 3'h0;
  assign v_4506_0 = v_4507_0 | v_4508_0;
  assign v_4507_0 = v_589_0 | v_601_0;
  assign v_4508_0 = v_607_0 | v_26_0;
  assign v_4509_0 = v_4510_0 | v_9765_0;
  assign v_4510_0 = v_4511_0 | v_9764_0;
  assign v_4511_0 = v_589_0 ? v_4512_0 : 3'h0;
  assign v_4513_0 = v_4514_0 | v_4515_0;
  assign v_4514_0 = v_589_0 | v_601_0;
  assign v_4515_0 = v_607_0 | v_26_0;
  assign v_4516_0 = v_4517_0 | v_9761_0;
  assign v_4517_0 = v_4518_0 | v_9760_0;
  assign v_4518_0 = v_589_0 ? v_4519_0 : 3'h0;
  assign v_4520_0 = v_4521_0 | v_4522_0;
  assign v_4521_0 = v_589_0 | v_601_0;
  assign v_4522_0 = v_607_0 | v_26_0;
  assign v_4523_0 = v_4524_0 | v_9757_0;
  assign v_4524_0 = v_4525_0 | v_9756_0;
  assign v_4525_0 = v_589_0 ? v_4526_0 : 3'h0;
  assign v_4527_0 = v_4528_0 | v_4529_0;
  assign v_4528_0 = v_589_0 | v_601_0;
  assign v_4529_0 = v_607_0 | v_26_0;
  assign v_4530_0 = v_4531_0 | v_9753_0;
  assign v_4531_0 = v_4532_0 | v_9752_0;
  assign v_4532_0 = v_589_0 ? v_4533_0 : 3'h0;
  assign v_4534_0 = v_4535_0 | v_4536_0;
  assign v_4535_0 = v_589_0 | v_601_0;
  assign v_4536_0 = v_607_0 | v_26_0;
  assign v_4537_0 = v_4538_0 | v_9749_0;
  assign v_4538_0 = v_4539_0 | v_9748_0;
  assign v_4539_0 = v_589_0 ? v_4540_0 : 3'h0;
  assign v_4541_0 = v_4542_0 | v_4543_0;
  assign v_4542_0 = v_589_0 | v_601_0;
  assign v_4543_0 = v_607_0 | v_26_0;
  assign v_4544_0 = v_4545_0 | v_9745_0;
  assign v_4545_0 = v_4546_0 | v_9744_0;
  assign v_4546_0 = v_589_0 ? v_4547_0 : 3'h0;
  assign v_4548_0 = v_4549_0 | v_4550_0;
  assign v_4549_0 = v_589_0 | v_601_0;
  assign v_4550_0 = v_607_0 | v_26_0;
  assign v_4551_0 = v_4552_0 | v_9741_0;
  assign v_4552_0 = v_4553_0 | v_9740_0;
  assign v_4553_0 = v_589_0 ? v_4554_0 : 3'h0;
  assign v_4555_0 = v_4556_0 | v_4557_0;
  assign v_4556_0 = v_589_0 | v_601_0;
  assign v_4557_0 = v_607_0 | v_26_0;
  assign v_4558_0 = v_4559_0 | v_9737_0;
  assign v_4559_0 = v_4560_0 | v_9736_0;
  assign v_4560_0 = v_589_0 ? v_4561_0 : 3'h0;
  assign v_4562_0 = v_4563_0 | v_4564_0;
  assign v_4563_0 = v_589_0 | v_601_0;
  assign v_4564_0 = v_607_0 | v_26_0;
  assign v_4565_0 = v_4566_0 | v_9733_0;
  assign v_4566_0 = v_4567_0 | v_9732_0;
  assign v_4567_0 = v_589_0 ? v_4568_0 : 3'h0;
  assign v_4569_0 = v_4570_0 | v_4571_0;
  assign v_4570_0 = v_589_0 | v_601_0;
  assign v_4571_0 = v_607_0 | v_26_0;
  assign v_4572_0 = v_4573_0 | v_9729_0;
  assign v_4573_0 = v_4574_0 | v_9728_0;
  assign v_4574_0 = v_589_0 ? v_4575_0 : 3'h0;
  assign v_4576_0 = v_4577_0 | v_4578_0;
  assign v_4577_0 = v_589_0 | v_601_0;
  assign v_4578_0 = v_607_0 | v_26_0;
  assign v_4579_0 = v_4580_0 | v_9725_0;
  assign v_4580_0 = v_4581_0 | v_9724_0;
  assign v_4581_0 = v_589_0 ? v_4582_0 : 3'h0;
  assign v_4583_0 = v_4584_0 | v_4585_0;
  assign v_4584_0 = v_589_0 | v_601_0;
  assign v_4585_0 = v_607_0 | v_26_0;
  assign v_4586_0 = v_4587_0 | v_9721_0;
  assign v_4587_0 = v_4588_0 | v_9720_0;
  assign v_4588_0 = v_589_0 ? v_4589_0 : 3'h0;
  assign v_4590_0 = v_4591_0 | v_4592_0;
  assign v_4591_0 = v_589_0 | v_601_0;
  assign v_4592_0 = v_607_0 | v_26_0;
  assign v_4593_0 = v_4594_0 | v_9717_0;
  assign v_4594_0 = v_4595_0 | v_9716_0;
  assign v_4595_0 = v_589_0 ? v_4596_0 : 3'h0;
  assign v_4597_0 = v_4598_0 | v_4599_0;
  assign v_4598_0 = v_589_0 | v_601_0;
  assign v_4599_0 = v_607_0 | v_26_0;
  assign v_4600_0 = v_4601_0 | v_9713_0;
  assign v_4601_0 = v_4602_0 | v_9712_0;
  assign v_4602_0 = v_589_0 ? v_4603_0 : 3'h0;
  assign v_4604_0 = v_4605_0 | v_4606_0;
  assign v_4605_0 = v_589_0 | v_601_0;
  assign v_4606_0 = v_607_0 | v_26_0;
  assign v_4607_0 = v_4608_0 | v_9709_0;
  assign v_4608_0 = v_4609_0 | v_9708_0;
  assign v_4609_0 = v_589_0 ? v_4610_0 : 3'h0;
  assign v_4611_0 = v_4612_0 | v_4613_0;
  assign v_4612_0 = v_589_0 | v_601_0;
  assign v_4613_0 = v_607_0 | v_26_0;
  assign v_4614_0 = v_4615_0 | v_9705_0;
  assign v_4615_0 = v_4616_0 | v_9704_0;
  assign v_4616_0 = v_589_0 ? v_4617_0 : 3'h0;
  assign v_4618_0 = v_4619_0 | v_4620_0;
  assign v_4619_0 = v_589_0 | v_601_0;
  assign v_4620_0 = v_607_0 | v_26_0;
  assign v_4621_0 = v_4622_0 | v_9701_0;
  assign v_4622_0 = v_4623_0 | v_9700_0;
  assign v_4623_0 = v_589_0 ? v_4624_0 : 3'h0;
  assign v_4625_0 = v_4626_0 | v_4627_0;
  assign v_4626_0 = v_589_0 | v_601_0;
  assign v_4627_0 = v_607_0 | v_26_0;
  assign v_4628_0 = v_4629_0 | v_9697_0;
  assign v_4629_0 = v_4630_0 | v_9696_0;
  assign v_4630_0 = v_589_0 ? v_4631_0 : 3'h0;
  assign v_4632_0 = v_4633_0 | v_4634_0;
  assign v_4633_0 = v_589_0 | v_601_0;
  assign v_4634_0 = v_607_0 | v_26_0;
  assign v_4635_0 = v_4636_0 | v_9693_0;
  assign v_4636_0 = v_4637_0 | v_9692_0;
  assign v_4637_0 = v_589_0 ? v_4638_0 : 3'h0;
  assign v_4639_0 = v_4640_0 | v_4641_0;
  assign v_4640_0 = v_589_0 | v_601_0;
  assign v_4641_0 = v_607_0 | v_26_0;
  assign v_4642_0 = v_4643_0 | v_9689_0;
  assign v_4643_0 = v_4644_0 | v_9688_0;
  assign v_4644_0 = v_589_0 ? v_4645_0 : 3'h0;
  assign v_4646_0 = v_4647_0 | v_4648_0;
  assign v_4647_0 = v_589_0 | v_601_0;
  assign v_4648_0 = v_607_0 | v_26_0;
  assign v_4649_0 = v_4650_0 | v_9685_0;
  assign v_4650_0 = v_4651_0 | v_9684_0;
  assign v_4651_0 = v_589_0 ? v_4652_0 : 3'h0;
  assign v_4653_0 = v_4654_0 | v_4655_0;
  assign v_4654_0 = v_589_0 | v_601_0;
  assign v_4655_0 = v_607_0 | v_26_0;
  assign v_4656_0 = v_4657_0 | v_9681_0;
  assign v_4657_0 = v_4658_0 | v_9680_0;
  assign v_4658_0 = v_589_0 ? v_4659_0 : 3'h0;
  assign v_4660_0 = v_4661_0 | v_4662_0;
  assign v_4661_0 = v_589_0 | v_601_0;
  assign v_4662_0 = v_607_0 | v_26_0;
  assign v_4663_0 = v_4664_0 | v_9677_0;
  assign v_4664_0 = v_4665_0 | v_9676_0;
  assign v_4665_0 = v_589_0 ? v_4666_0 : 3'h0;
  assign v_4667_0 = v_4668_0 | v_4669_0;
  assign v_4668_0 = v_589_0 | v_601_0;
  assign v_4669_0 = v_607_0 | v_26_0;
  assign v_4670_0 = v_4671_0 | v_9673_0;
  assign v_4671_0 = v_4672_0 | v_9672_0;
  assign v_4672_0 = v_589_0 ? v_4673_0 : 3'h0;
  assign v_4674_0 = v_4675_0 | v_4676_0;
  assign v_4675_0 = v_589_0 | v_601_0;
  assign v_4676_0 = v_607_0 | v_26_0;
  assign v_4677_0 = v_4678_0 | v_9669_0;
  assign v_4678_0 = v_4679_0 | v_9668_0;
  assign v_4679_0 = v_589_0 ? v_4680_0 : 3'h0;
  assign v_4681_0 = v_4682_0 | v_4683_0;
  assign v_4682_0 = v_589_0 | v_601_0;
  assign v_4683_0 = v_607_0 | v_26_0;
  assign v_4684_0 = v_4685_0 | v_9665_0;
  assign v_4685_0 = v_4686_0 | v_9664_0;
  assign v_4686_0 = v_589_0 ? v_4687_0 : 3'h0;
  assign v_4688_0 = v_4689_0 | v_4690_0;
  assign v_4689_0 = v_589_0 | v_601_0;
  assign v_4690_0 = v_607_0 | v_26_0;
  assign v_4691_0 = v_4692_0 | v_9661_0;
  assign v_4692_0 = v_4693_0 | v_9660_0;
  assign v_4693_0 = v_589_0 ? v_4694_0 : 3'h0;
  assign v_4695_0 = v_4696_0 | v_4697_0;
  assign v_4696_0 = v_589_0 | v_601_0;
  assign v_4697_0 = v_607_0 | v_26_0;
  assign v_4698_0 = v_4699_0 | v_9657_0;
  assign v_4699_0 = v_4700_0 | v_9656_0;
  assign v_4700_0 = v_589_0 ? v_4701_0 : 3'h0;
  assign v_4702_0 = v_4703_0 | v_4704_0;
  assign v_4703_0 = v_589_0 | v_601_0;
  assign v_4704_0 = v_607_0 | v_26_0;
  assign v_4705_0 = v_4706_0 | v_9653_0;
  assign v_4706_0 = v_4707_0 | v_9652_0;
  assign v_4707_0 = v_589_0 ? v_4708_0 : 3'h0;
  assign v_4709_0 = v_4710_0 | v_4711_0;
  assign v_4710_0 = v_589_0 | v_601_0;
  assign v_4711_0 = v_607_0 | v_26_0;
  assign v_4712_0 = v_4713_0 | v_9649_0;
  assign v_4713_0 = v_4714_0 | v_9648_0;
  assign v_4714_0 = v_589_0 ? v_4715_0 : 3'h0;
  assign v_4716_0 = v_4717_0 | v_4718_0;
  assign v_4717_0 = v_589_0 | v_601_0;
  assign v_4718_0 = v_607_0 | v_26_0;
  assign v_4719_0 = v_4720_0 | v_9645_0;
  assign v_4720_0 = v_4721_0 | v_9644_0;
  assign v_4721_0 = v_589_0 ? v_4722_0 : 3'h0;
  assign v_4723_0 = v_4724_0 | v_4725_0;
  assign v_4724_0 = v_589_0 | v_601_0;
  assign v_4725_0 = v_607_0 | v_26_0;
  assign v_4726_0 = v_4727_0 | v_9641_0;
  assign v_4727_0 = v_4728_0 | v_9640_0;
  assign v_4728_0 = v_589_0 ? v_4729_0 : 3'h0;
  assign v_4730_0 = v_4731_0 | v_4732_0;
  assign v_4731_0 = v_589_0 | v_601_0;
  assign v_4732_0 = v_607_0 | v_26_0;
  assign v_4733_0 = v_4734_0 | v_9637_0;
  assign v_4734_0 = v_4735_0 | v_9636_0;
  assign v_4735_0 = v_589_0 ? v_4736_0 : 3'h0;
  assign v_4737_0 = v_4738_0 | v_4739_0;
  assign v_4738_0 = v_589_0 | v_601_0;
  assign v_4739_0 = v_607_0 | v_26_0;
  assign v_4740_0 = v_4741_0 | v_9633_0;
  assign v_4741_0 = v_4742_0 | v_9632_0;
  assign v_4742_0 = v_589_0 ? v_4743_0 : 3'h0;
  assign v_4744_0 = v_4745_0 | v_4746_0;
  assign v_4745_0 = v_589_0 | v_601_0;
  assign v_4746_0 = v_607_0 | v_26_0;
  assign v_4747_0 = v_4748_0 | v_9629_0;
  assign v_4748_0 = v_4749_0 | v_9628_0;
  assign v_4749_0 = v_589_0 ? v_4750_0 : 3'h0;
  assign v_4751_0 = v_4752_0 | v_4753_0;
  assign v_4752_0 = v_589_0 | v_601_0;
  assign v_4753_0 = v_607_0 | v_26_0;
  assign v_4754_0 = v_4755_0 | v_9625_0;
  assign v_4755_0 = v_4756_0 | v_9624_0;
  assign v_4756_0 = v_589_0 ? v_4757_0 : 3'h0;
  assign v_4758_0 = v_4759_0 | v_4760_0;
  assign v_4759_0 = v_589_0 | v_601_0;
  assign v_4760_0 = v_607_0 | v_26_0;
  assign v_4761_0 = v_4762_0 | v_9621_0;
  assign v_4762_0 = v_4763_0 | v_9620_0;
  assign v_4763_0 = v_589_0 ? v_4764_0 : 3'h0;
  assign v_4765_0 = v_4766_0 | v_4767_0;
  assign v_4766_0 = v_589_0 | v_601_0;
  assign v_4767_0 = v_607_0 | v_26_0;
  assign v_4768_0 = v_4769_0 | v_9617_0;
  assign v_4769_0 = v_4770_0 | v_9616_0;
  assign v_4770_0 = v_589_0 ? v_4771_0 : 3'h0;
  assign v_4772_0 = v_4773_0 | v_4774_0;
  assign v_4773_0 = v_589_0 | v_601_0;
  assign v_4774_0 = v_607_0 | v_26_0;
  assign v_4775_0 = v_4776_0 | v_9613_0;
  assign v_4776_0 = v_4777_0 | v_9612_0;
  assign v_4777_0 = v_589_0 ? v_4778_0 : 3'h0;
  assign v_4779_0 = v_4780_0 | v_4781_0;
  assign v_4780_0 = v_589_0 | v_601_0;
  assign v_4781_0 = v_607_0 | v_26_0;
  assign v_4782_0 = v_4783_0 | v_9609_0;
  assign v_4783_0 = v_4784_0 | v_9608_0;
  assign v_4784_0 = v_589_0 ? v_4785_0 : 3'h0;
  assign v_4786_0 = v_4787_0 | v_4788_0;
  assign v_4787_0 = v_589_0 | v_601_0;
  assign v_4788_0 = v_607_0 | v_26_0;
  assign v_4789_0 = v_4790_0 | v_9605_0;
  assign v_4790_0 = v_4791_0 | v_9604_0;
  assign v_4791_0 = v_589_0 ? v_4792_0 : 3'h0;
  assign v_4793_0 = v_4794_0 | v_4795_0;
  assign v_4794_0 = v_589_0 | v_601_0;
  assign v_4795_0 = v_607_0 | v_26_0;
  assign v_4796_0 = v_4797_0 | v_9601_0;
  assign v_4797_0 = v_4798_0 | v_9600_0;
  assign v_4798_0 = v_589_0 ? v_4799_0 : 3'h0;
  assign v_4800_0 = v_4801_0 | v_4802_0;
  assign v_4801_0 = v_589_0 | v_601_0;
  assign v_4802_0 = v_607_0 | v_26_0;
  assign v_4803_0 = v_4804_0 | v_9597_0;
  assign v_4804_0 = v_4805_0 | v_9596_0;
  assign v_4805_0 = v_589_0 ? v_4806_0 : 3'h0;
  assign v_4807_0 = v_4808_0 | v_4809_0;
  assign v_4808_0 = v_589_0 | v_601_0;
  assign v_4809_0 = v_607_0 | v_26_0;
  assign v_4810_0 = v_4811_0 | v_9593_0;
  assign v_4811_0 = v_4812_0 | v_9592_0;
  assign v_4812_0 = v_589_0 ? v_4813_0 : 3'h0;
  assign v_4814_0 = v_4815_0 | v_4816_0;
  assign v_4815_0 = v_589_0 | v_601_0;
  assign v_4816_0 = v_607_0 | v_26_0;
  assign v_4817_0 = v_4818_0 | v_9589_0;
  assign v_4818_0 = v_4819_0 | v_9588_0;
  assign v_4819_0 = v_589_0 ? v_4820_0 : 3'h0;
  assign v_4821_0 = v_4822_0 | v_4823_0;
  assign v_4822_0 = v_589_0 | v_601_0;
  assign v_4823_0 = v_607_0 | v_26_0;
  assign v_4824_0 = v_4825_0 | v_9585_0;
  assign v_4825_0 = v_4826_0 | v_9584_0;
  assign v_4826_0 = v_589_0 ? v_4827_0 : 3'h0;
  assign v_4828_0 = v_4829_0 | v_4830_0;
  assign v_4829_0 = v_589_0 | v_601_0;
  assign v_4830_0 = v_607_0 | v_26_0;
  assign v_4831_0 = v_4832_0 | v_9581_0;
  assign v_4832_0 = v_4833_0 | v_9580_0;
  assign v_4833_0 = v_589_0 ? v_4834_0 : 3'h0;
  assign v_4835_0 = v_4836_0 | v_4837_0;
  assign v_4836_0 = v_589_0 | v_601_0;
  assign v_4837_0 = v_607_0 | v_26_0;
  assign v_4838_0 = v_4839_0 | v_9577_0;
  assign v_4839_0 = v_4840_0 | v_9576_0;
  assign v_4840_0 = v_589_0 ? v_4841_0 : 3'h0;
  assign v_4842_0 = v_4843_0 | v_4844_0;
  assign v_4843_0 = v_589_0 | v_601_0;
  assign v_4844_0 = v_607_0 | v_26_0;
  assign v_4845_0 = v_4846_0 | v_9573_0;
  assign v_4846_0 = v_4847_0 | v_9572_0;
  assign v_4847_0 = v_589_0 ? v_4848_0 : 3'h0;
  assign v_4849_0 = v_4850_0 | v_4851_0;
  assign v_4850_0 = v_589_0 | v_601_0;
  assign v_4851_0 = v_607_0 | v_26_0;
  assign v_4852_0 = v_4853_0 | v_9569_0;
  assign v_4853_0 = v_4854_0 | v_9568_0;
  assign v_4854_0 = v_589_0 ? v_4855_0 : 3'h0;
  assign v_4856_0 = v_4857_0 | v_4858_0;
  assign v_4857_0 = v_589_0 | v_601_0;
  assign v_4858_0 = v_607_0 | v_26_0;
  assign v_4859_0 = v_4860_0 | v_9565_0;
  assign v_4860_0 = v_4861_0 | v_9564_0;
  assign v_4861_0 = v_589_0 ? v_4862_0 : 3'h0;
  assign v_4863_0 = v_4864_0 | v_4865_0;
  assign v_4864_0 = v_589_0 | v_601_0;
  assign v_4865_0 = v_607_0 | v_26_0;
  assign v_4866_0 = v_4867_0 | v_9561_0;
  assign v_4867_0 = v_4868_0 | v_9560_0;
  assign v_4868_0 = v_589_0 ? v_4869_0 : 3'h0;
  assign v_4870_0 = v_4871_0 | v_4872_0;
  assign v_4871_0 = v_589_0 | v_601_0;
  assign v_4872_0 = v_607_0 | v_26_0;
  assign v_4873_0 = v_4874_0 | v_9557_0;
  assign v_4874_0 = v_4875_0 | v_9556_0;
  assign v_4875_0 = v_589_0 ? v_4876_0 : 3'h0;
  assign v_4877_0 = v_4878_0 | v_4879_0;
  assign v_4878_0 = v_589_0 | v_601_0;
  assign v_4879_0 = v_607_0 | v_26_0;
  assign v_4880_0 = v_4881_0 | v_9553_0;
  assign v_4881_0 = v_4882_0 | v_9552_0;
  assign v_4882_0 = v_589_0 ? v_4883_0 : 3'h0;
  assign v_4884_0 = v_4885_0 | v_4886_0;
  assign v_4885_0 = v_589_0 | v_601_0;
  assign v_4886_0 = v_607_0 | v_26_0;
  assign v_4887_0 = v_4888_0 | v_9549_0;
  assign v_4888_0 = v_4889_0 | v_9548_0;
  assign v_4889_0 = v_589_0 ? v_4890_0 : 3'h0;
  assign v_4891_0 = v_4892_0 | v_4893_0;
  assign v_4892_0 = v_589_0 | v_601_0;
  assign v_4893_0 = v_607_0 | v_26_0;
  assign v_4894_0 = v_4895_0 | v_9545_0;
  assign v_4895_0 = v_4896_0 | v_9544_0;
  assign v_4896_0 = v_589_0 ? v_4897_0 : 3'h0;
  assign v_4898_0 = v_4899_0 | v_4900_0;
  assign v_4899_0 = v_589_0 | v_601_0;
  assign v_4900_0 = v_607_0 | v_26_0;
  assign v_4901_0 = v_4902_0 | v_9541_0;
  assign v_4902_0 = v_4903_0 | v_9540_0;
  assign v_4903_0 = v_589_0 ? v_4904_0 : 3'h0;
  assign v_4905_0 = v_4906_0 | v_4907_0;
  assign v_4906_0 = v_589_0 | v_601_0;
  assign v_4907_0 = v_607_0 | v_26_0;
  assign v_4908_0 = v_4909_0 | v_9537_0;
  assign v_4909_0 = v_4910_0 | v_9536_0;
  assign v_4910_0 = v_589_0 ? v_4911_0 : 3'h0;
  assign v_4912_0 = v_4913_0 | v_4914_0;
  assign v_4913_0 = v_589_0 | v_601_0;
  assign v_4914_0 = v_607_0 | v_26_0;
  assign v_4915_0 = v_4916_0 | v_9533_0;
  assign v_4916_0 = v_4917_0 | v_9532_0;
  assign v_4917_0 = v_589_0 ? v_4918_0 : 3'h0;
  assign v_4919_0 = v_4920_0 | v_4921_0;
  assign v_4920_0 = v_589_0 | v_601_0;
  assign v_4921_0 = v_607_0 | v_26_0;
  assign v_4922_0 = v_4923_0 | v_9529_0;
  assign v_4923_0 = v_4924_0 | v_9528_0;
  assign v_4924_0 = v_589_0 ? v_4925_0 : 3'h0;
  assign v_4926_0 = v_4927_0 | v_4928_0;
  assign v_4927_0 = v_589_0 | v_601_0;
  assign v_4928_0 = v_607_0 | v_26_0;
  assign v_4929_0 = v_4930_0 | v_9525_0;
  assign v_4930_0 = v_4931_0 | v_9524_0;
  assign v_4931_0 = v_589_0 ? v_4932_0 : 3'h0;
  assign v_4933_0 = v_4934_0 | v_4935_0;
  assign v_4934_0 = v_589_0 | v_601_0;
  assign v_4935_0 = v_607_0 | v_26_0;
  assign v_4936_0 = v_4937_0 | v_9521_0;
  assign v_4937_0 = v_4938_0 | v_9520_0;
  assign v_4938_0 = v_589_0 ? v_4939_0 : 3'h0;
  assign v_4940_0 = v_4941_0 | v_4942_0;
  assign v_4941_0 = v_589_0 | v_601_0;
  assign v_4942_0 = v_607_0 | v_26_0;
  assign v_4943_0 = v_4944_0 | v_9517_0;
  assign v_4944_0 = v_4945_0 | v_9516_0;
  assign v_4945_0 = v_589_0 ? v_4946_0 : 3'h0;
  assign v_4947_0 = v_4948_0 | v_4949_0;
  assign v_4948_0 = v_589_0 | v_601_0;
  assign v_4949_0 = v_607_0 | v_26_0;
  assign v_4950_0 = v_4951_0 | v_9513_0;
  assign v_4951_0 = v_4952_0 | v_9512_0;
  assign v_4952_0 = v_589_0 ? v_4953_0 : 3'h0;
  assign v_4954_0 = v_4955_0 | v_4956_0;
  assign v_4955_0 = v_589_0 | v_601_0;
  assign v_4956_0 = v_607_0 | v_26_0;
  assign v_4957_0 = v_4958_0 | v_9509_0;
  assign v_4958_0 = v_4959_0 | v_9508_0;
  assign v_4959_0 = v_589_0 ? v_4960_0 : 3'h0;
  assign v_4961_0 = v_4962_0 | v_4963_0;
  assign v_4962_0 = v_589_0 | v_601_0;
  assign v_4963_0 = v_607_0 | v_26_0;
  assign v_4964_0 = v_4965_0 | v_9505_0;
  assign v_4965_0 = v_4966_0 | v_9504_0;
  assign v_4966_0 = v_589_0 ? v_4967_0 : 3'h0;
  assign v_4968_0 = v_4969_0 | v_4970_0;
  assign v_4969_0 = v_589_0 | v_601_0;
  assign v_4970_0 = v_607_0 | v_26_0;
  assign v_4971_0 = v_4972_0 | v_9501_0;
  assign v_4972_0 = v_4973_0 | v_9500_0;
  assign v_4973_0 = v_589_0 ? v_4974_0 : 3'h0;
  assign v_4975_0 = v_4976_0 | v_4977_0;
  assign v_4976_0 = v_589_0 | v_601_0;
  assign v_4977_0 = v_607_0 | v_26_0;
  assign v_4978_0 = v_4979_0 | v_9497_0;
  assign v_4979_0 = v_4980_0 | v_9496_0;
  assign v_4980_0 = v_589_0 ? v_4981_0 : 3'h0;
  assign v_4982_0 = v_4983_0 | v_4984_0;
  assign v_4983_0 = v_589_0 | v_601_0;
  assign v_4984_0 = v_607_0 | v_26_0;
  assign v_4985_0 = v_4986_0 | v_9493_0;
  assign v_4986_0 = v_4987_0 | v_9492_0;
  assign v_4987_0 = v_589_0 ? v_4988_0 : 3'h0;
  assign v_4989_0 = v_4990_0 | v_4991_0;
  assign v_4990_0 = v_589_0 | v_601_0;
  assign v_4991_0 = v_607_0 | v_26_0;
  assign v_4992_0 = v_4993_0 | v_9489_0;
  assign v_4993_0 = v_4994_0 | v_9488_0;
  assign v_4994_0 = v_589_0 ? v_4995_0 : 3'h0;
  assign v_4996_0 = v_4997_0 | v_4998_0;
  assign v_4997_0 = v_589_0 | v_601_0;
  assign v_4998_0 = v_607_0 | v_26_0;
  assign v_4999_0 = v_5000_0 | v_9485_0;
  assign v_5000_0 = v_5001_0 | v_9484_0;
  assign v_5001_0 = v_589_0 ? v_5002_0 : 3'h0;
  assign v_5003_0 = v_5004_0 | v_5005_0;
  assign v_5004_0 = v_589_0 | v_601_0;
  assign v_5005_0 = v_607_0 | v_26_0;
  assign v_5006_0 = v_5007_0 | v_9481_0;
  assign v_5007_0 = v_5008_0 | v_9480_0;
  assign v_5008_0 = v_589_0 ? v_5009_0 : 3'h0;
  assign v_5010_0 = v_5011_0 | v_5012_0;
  assign v_5011_0 = v_589_0 | v_601_0;
  assign v_5012_0 = v_607_0 | v_26_0;
  assign v_5013_0 = v_5014_0 | v_9477_0;
  assign v_5014_0 = v_5015_0 | v_9476_0;
  assign v_5015_0 = v_589_0 ? v_5016_0 : 3'h0;
  assign v_5017_0 = v_5018_0 | v_5019_0;
  assign v_5018_0 = v_589_0 | v_601_0;
  assign v_5019_0 = v_607_0 | v_26_0;
  assign v_5020_0 = v_5021_0 | v_9473_0;
  assign v_5021_0 = v_5022_0 | v_9472_0;
  assign v_5022_0 = v_589_0 ? v_5023_0 : 3'h0;
  assign v_5024_0 = v_5025_0 | v_5026_0;
  assign v_5025_0 = v_589_0 | v_601_0;
  assign v_5026_0 = v_607_0 | v_26_0;
  assign v_5027_0 = v_5028_0 | v_9469_0;
  assign v_5028_0 = v_5029_0 | v_9468_0;
  assign v_5029_0 = v_589_0 ? v_5030_0 : 3'h0;
  assign v_5031_0 = v_5032_0 | v_5033_0;
  assign v_5032_0 = v_589_0 | v_601_0;
  assign v_5033_0 = v_607_0 | v_26_0;
  assign v_5034_0 = v_5035_0 | v_9465_0;
  assign v_5035_0 = v_5036_0 | v_9464_0;
  assign v_5036_0 = v_589_0 ? v_5037_0 : 3'h0;
  assign v_5038_0 = v_5039_0 | v_5040_0;
  assign v_5039_0 = v_589_0 | v_601_0;
  assign v_5040_0 = v_607_0 | v_26_0;
  assign v_5041_0 = v_5042_0 | v_9461_0;
  assign v_5042_0 = v_5043_0 | v_9460_0;
  assign v_5043_0 = v_589_0 ? v_5044_0 : 3'h0;
  assign v_5045_0 = v_5046_0 | v_5047_0;
  assign v_5046_0 = v_589_0 | v_601_0;
  assign v_5047_0 = v_607_0 | v_26_0;
  assign v_5048_0 = v_5049_0 | v_9457_0;
  assign v_5049_0 = v_5050_0 | v_9456_0;
  assign v_5050_0 = v_589_0 ? v_5051_0 : 3'h0;
  assign v_5052_0 = v_5053_0 | v_5054_0;
  assign v_5053_0 = v_589_0 | v_601_0;
  assign v_5054_0 = v_607_0 | v_26_0;
  assign v_5055_0 = v_5056_0 | v_9453_0;
  assign v_5056_0 = v_5057_0 | v_9452_0;
  assign v_5057_0 = v_589_0 ? v_5058_0 : 3'h0;
  assign v_5059_0 = v_5060_0 | v_5061_0;
  assign v_5060_0 = v_589_0 | v_601_0;
  assign v_5061_0 = v_607_0 | v_26_0;
  assign v_5062_0 = v_5063_0 | v_9449_0;
  assign v_5063_0 = v_5064_0 | v_9448_0;
  assign v_5064_0 = v_589_0 ? v_5065_0 : 3'h0;
  assign v_5066_0 = v_5067_0 | v_5068_0;
  assign v_5067_0 = v_589_0 | v_601_0;
  assign v_5068_0 = v_607_0 | v_26_0;
  assign v_5069_0 = v_5070_0 | v_9445_0;
  assign v_5070_0 = v_5071_0 | v_9444_0;
  assign v_5071_0 = v_589_0 ? v_5072_0 : 3'h0;
  assign v_5073_0 = v_5074_0 | v_5075_0;
  assign v_5074_0 = v_589_0 | v_601_0;
  assign v_5075_0 = v_607_0 | v_26_0;
  assign v_5076_0 = v_5077_0 | v_9441_0;
  assign v_5077_0 = v_5078_0 | v_9440_0;
  assign v_5078_0 = v_589_0 ? v_5079_0 : 3'h0;
  assign v_5080_0 = v_5081_0 | v_5082_0;
  assign v_5081_0 = v_589_0 | v_601_0;
  assign v_5082_0 = v_607_0 | v_26_0;
  assign v_5083_0 = v_5084_0 | v_9437_0;
  assign v_5084_0 = v_5085_0 | v_9436_0;
  assign v_5085_0 = v_589_0 ? v_5086_0 : 3'h0;
  assign v_5087_0 = v_5088_0 | v_5089_0;
  assign v_5088_0 = v_589_0 | v_601_0;
  assign v_5089_0 = v_607_0 | v_26_0;
  assign v_5090_0 = v_5091_0 | v_9433_0;
  assign v_5091_0 = v_5092_0 | v_9432_0;
  assign v_5092_0 = v_589_0 ? v_5093_0 : 3'h0;
  assign v_5094_0 = v_5095_0 | v_5096_0;
  assign v_5095_0 = v_589_0 | v_601_0;
  assign v_5096_0 = v_607_0 | v_26_0;
  assign v_5097_0 = v_5098_0 | v_9429_0;
  assign v_5098_0 = v_5099_0 | v_9428_0;
  assign v_5099_0 = v_589_0 ? v_5100_0 : 3'h0;
  assign v_5101_0 = v_5102_0 | v_5103_0;
  assign v_5102_0 = v_589_0 | v_601_0;
  assign v_5103_0 = v_607_0 | v_26_0;
  assign v_5104_0 = v_5105_0 | v_9425_0;
  assign v_5105_0 = v_5106_0 | v_9424_0;
  assign v_5106_0 = v_589_0 ? v_5107_0 : 3'h0;
  assign v_5108_0 = v_5109_0 | v_5110_0;
  assign v_5109_0 = v_589_0 | v_601_0;
  assign v_5110_0 = v_607_0 | v_26_0;
  assign v_5111_0 = v_5112_0 | v_9421_0;
  assign v_5112_0 = v_5113_0 | v_9420_0;
  assign v_5113_0 = v_589_0 ? v_5114_0 : 3'h0;
  assign v_5115_0 = v_5116_0 | v_5117_0;
  assign v_5116_0 = v_589_0 | v_601_0;
  assign v_5117_0 = v_607_0 | v_26_0;
  assign v_5118_0 = v_5119_0 | v_9417_0;
  assign v_5119_0 = v_5120_0 | v_9416_0;
  assign v_5120_0 = v_589_0 ? v_5121_0 : 3'h0;
  assign v_5122_0 = v_5123_0 | v_5124_0;
  assign v_5123_0 = v_589_0 | v_601_0;
  assign v_5124_0 = v_607_0 | v_26_0;
  assign v_5125_0 = v_5126_0 | v_9413_0;
  assign v_5126_0 = v_5127_0 | v_9412_0;
  assign v_5127_0 = v_589_0 ? v_5128_0 : 3'h0;
  assign v_5129_0 = v_5130_0 | v_5131_0;
  assign v_5130_0 = v_589_0 | v_601_0;
  assign v_5131_0 = v_607_0 | v_26_0;
  assign v_5132_0 = v_5133_0 | v_9409_0;
  assign v_5133_0 = v_5134_0 | v_9408_0;
  assign v_5134_0 = v_589_0 ? v_5135_0 : 3'h0;
  assign v_5136_0 = v_5137_0 | v_5138_0;
  assign v_5137_0 = v_589_0 | v_601_0;
  assign v_5138_0 = v_607_0 | v_26_0;
  assign v_5139_0 = v_5140_0 | v_9405_0;
  assign v_5140_0 = v_5141_0 | v_9404_0;
  assign v_5141_0 = v_589_0 ? v_5142_0 : 3'h0;
  assign v_5143_0 = v_5144_0 | v_5145_0;
  assign v_5144_0 = v_589_0 | v_601_0;
  assign v_5145_0 = v_607_0 | v_26_0;
  assign v_5146_0 = v_5147_0 | v_9401_0;
  assign v_5147_0 = v_5148_0 | v_9400_0;
  assign v_5148_0 = v_589_0 ? v_5149_0 : 3'h0;
  assign v_5150_0 = v_5151_0 | v_5152_0;
  assign v_5151_0 = v_589_0 | v_601_0;
  assign v_5152_0 = v_607_0 | v_26_0;
  assign v_5153_0 = v_5154_0 | v_9397_0;
  assign v_5154_0 = v_5155_0 | v_9396_0;
  assign v_5155_0 = v_589_0 ? v_5156_0 : 3'h0;
  assign v_5157_0 = v_5158_0 | v_5159_0;
  assign v_5158_0 = v_589_0 | v_601_0;
  assign v_5159_0 = v_607_0 | v_26_0;
  assign v_5160_0 = v_5161_0 | v_9393_0;
  assign v_5161_0 = v_5162_0 | v_9392_0;
  assign v_5162_0 = v_589_0 ? v_5163_0 : 3'h0;
  assign v_5164_0 = v_5165_0 | v_5166_0;
  assign v_5165_0 = v_589_0 | v_601_0;
  assign v_5166_0 = v_607_0 | v_26_0;
  assign v_5167_0 = v_5168_0 | v_9389_0;
  assign v_5168_0 = v_5169_0 | v_9388_0;
  assign v_5169_0 = v_589_0 ? v_5170_0 : 3'h0;
  assign v_5171_0 = v_5172_0 | v_5173_0;
  assign v_5172_0 = v_589_0 | v_601_0;
  assign v_5173_0 = v_607_0 | v_26_0;
  assign v_5174_0 = v_5175_0 | v_9385_0;
  assign v_5175_0 = v_5176_0 | v_9384_0;
  assign v_5176_0 = v_589_0 ? v_5177_0 : 3'h0;
  assign v_5178_0 = v_5179_0 | v_5180_0;
  assign v_5179_0 = v_589_0 | v_601_0;
  assign v_5180_0 = v_607_0 | v_26_0;
  assign v_5181_0 = v_5182_0 | v_9381_0;
  assign v_5182_0 = v_5183_0 | v_9380_0;
  assign v_5183_0 = v_589_0 ? v_5184_0 : 3'h0;
  assign v_5185_0 = v_5186_0 | v_5187_0;
  assign v_5186_0 = v_589_0 | v_601_0;
  assign v_5187_0 = v_607_0 | v_26_0;
  assign v_5188_0 = v_5189_0 | v_9377_0;
  assign v_5189_0 = v_5190_0 | v_9376_0;
  assign v_5190_0 = v_589_0 ? v_5191_0 : 3'h0;
  assign v_5192_0 = v_5193_0 | v_5194_0;
  assign v_5193_0 = v_589_0 | v_601_0;
  assign v_5194_0 = v_607_0 | v_26_0;
  assign v_5195_0 = v_5196_0 | v_9373_0;
  assign v_5196_0 = v_5197_0 | v_9372_0;
  assign v_5197_0 = v_589_0 ? v_5198_0 : 3'h0;
  assign v_5199_0 = v_5200_0 | v_5201_0;
  assign v_5200_0 = v_589_0 | v_601_0;
  assign v_5201_0 = v_607_0 | v_26_0;
  assign v_5202_0 = v_5203_0 | v_9369_0;
  assign v_5203_0 = v_5204_0 | v_9368_0;
  assign v_5204_0 = v_589_0 ? v_5205_0 : 3'h0;
  assign v_5206_0 = v_5207_0 | v_5208_0;
  assign v_5207_0 = v_589_0 | v_601_0;
  assign v_5208_0 = v_607_0 | v_26_0;
  assign v_5209_0 = v_5210_0 | v_9365_0;
  assign v_5210_0 = v_5211_0 | v_9364_0;
  assign v_5211_0 = v_589_0 ? v_5212_0 : 3'h0;
  assign v_5213_0 = v_5214_0 | v_5215_0;
  assign v_5214_0 = v_589_0 | v_601_0;
  assign v_5215_0 = v_607_0 | v_26_0;
  assign v_5216_0 = v_5217_0 | v_9361_0;
  assign v_5217_0 = v_5218_0 | v_9360_0;
  assign v_5218_0 = v_589_0 ? v_5219_0 : 3'h0;
  assign v_5220_0 = v_5221_0 | v_5222_0;
  assign v_5221_0 = v_589_0 | v_601_0;
  assign v_5222_0 = v_607_0 | v_26_0;
  assign v_5223_0 = v_5224_0 | v_9357_0;
  assign v_5224_0 = v_5225_0 | v_9356_0;
  assign v_5225_0 = v_589_0 ? v_5226_0 : 3'h0;
  assign v_5227_0 = v_5228_0 | v_5229_0;
  assign v_5228_0 = v_589_0 | v_601_0;
  assign v_5229_0 = v_607_0 | v_26_0;
  assign v_5230_0 = v_5231_0 | v_9353_0;
  assign v_5231_0 = v_5232_0 | v_9352_0;
  assign v_5232_0 = v_589_0 ? v_5233_0 : 3'h0;
  assign v_5234_0 = v_5235_0 | v_5236_0;
  assign v_5235_0 = v_589_0 | v_601_0;
  assign v_5236_0 = v_607_0 | v_26_0;
  assign v_5237_0 = v_5238_0 | v_9349_0;
  assign v_5238_0 = v_5239_0 | v_9348_0;
  assign v_5239_0 = v_589_0 ? v_5240_0 : 3'h0;
  assign v_5241_0 = v_5242_0 | v_5243_0;
  assign v_5242_0 = v_589_0 | v_601_0;
  assign v_5243_0 = v_607_0 | v_26_0;
  assign v_5244_0 = v_5245_0 | v_9345_0;
  assign v_5245_0 = v_5246_0 | v_9344_0;
  assign v_5246_0 = v_589_0 ? v_5247_0 : 3'h0;
  assign v_5248_0 = v_5249_0 | v_5250_0;
  assign v_5249_0 = v_589_0 | v_601_0;
  assign v_5250_0 = v_607_0 | v_26_0;
  assign v_5251_0 = v_5252_0 | v_9341_0;
  assign v_5252_0 = v_5253_0 | v_9340_0;
  assign v_5253_0 = v_589_0 ? v_5254_0 : 3'h0;
  assign v_5255_0 = v_5256_0 | v_5257_0;
  assign v_5256_0 = v_589_0 | v_601_0;
  assign v_5257_0 = v_607_0 | v_26_0;
  assign v_5258_0 = v_5259_0 | v_9337_0;
  assign v_5259_0 = v_5260_0 | v_9336_0;
  assign v_5260_0 = v_589_0 ? v_5261_0 : 3'h0;
  assign v_5262_0 = v_5263_0 | v_5264_0;
  assign v_5263_0 = v_589_0 | v_601_0;
  assign v_5264_0 = v_607_0 | v_26_0;
  assign v_5265_0 = v_5266_0 | v_9333_0;
  assign v_5266_0 = v_5267_0 | v_9332_0;
  assign v_5267_0 = v_589_0 ? v_5268_0 : 3'h0;
  assign v_5269_0 = v_5270_0 | v_5271_0;
  assign v_5270_0 = v_589_0 | v_601_0;
  assign v_5271_0 = v_607_0 | v_26_0;
  assign v_5272_0 = v_5273_0 | v_9329_0;
  assign v_5273_0 = v_5274_0 | v_9328_0;
  assign v_5274_0 = v_589_0 ? v_5275_0 : 3'h0;
  assign v_5276_0 = v_5277_0 | v_5278_0;
  assign v_5277_0 = v_589_0 | v_601_0;
  assign v_5278_0 = v_607_0 | v_26_0;
  assign v_5279_0 = v_5280_0 | v_9325_0;
  assign v_5280_0 = v_5281_0 | v_9324_0;
  assign v_5281_0 = v_589_0 ? v_5282_0 : 3'h0;
  assign v_5283_0 = v_5284_0 | v_5285_0;
  assign v_5284_0 = v_589_0 | v_601_0;
  assign v_5285_0 = v_607_0 | v_26_0;
  assign v_5286_0 = v_5287_0 | v_9321_0;
  assign v_5287_0 = v_5288_0 | v_9320_0;
  assign v_5288_0 = v_589_0 ? v_5289_0 : 3'h0;
  assign v_5290_0 = v_5291_0 | v_5292_0;
  assign v_5291_0 = v_589_0 | v_601_0;
  assign v_5292_0 = v_607_0 | v_26_0;
  assign v_5293_0 = v_5294_0 | v_9317_0;
  assign v_5294_0 = v_5295_0 | v_9316_0;
  assign v_5295_0 = v_589_0 ? v_5296_0 : 3'h0;
  assign v_5297_0 = v_5298_0 | v_5299_0;
  assign v_5298_0 = v_589_0 | v_601_0;
  assign v_5299_0 = v_607_0 | v_26_0;
  assign v_5300_0 = v_5301_0 | v_9313_0;
  assign v_5301_0 = v_5302_0 | v_9312_0;
  assign v_5302_0 = v_589_0 ? v_5303_0 : 3'h0;
  assign v_5304_0 = v_5305_0 | v_5306_0;
  assign v_5305_0 = v_589_0 | v_601_0;
  assign v_5306_0 = v_607_0 | v_26_0;
  assign v_5307_0 = v_5308_0 | v_9309_0;
  assign v_5308_0 = v_5309_0 | v_9308_0;
  assign v_5309_0 = v_589_0 ? v_5310_0 : 3'h0;
  assign v_5311_0 = v_5312_0 | v_5313_0;
  assign v_5312_0 = v_589_0 | v_601_0;
  assign v_5313_0 = v_607_0 | v_26_0;
  assign v_5314_0 = v_5315_0 | v_9305_0;
  assign v_5315_0 = v_5316_0 | v_9304_0;
  assign v_5316_0 = v_589_0 ? v_5317_0 : 3'h0;
  assign v_5318_0 = v_5319_0 | v_5320_0;
  assign v_5319_0 = v_589_0 | v_601_0;
  assign v_5320_0 = v_607_0 | v_26_0;
  assign v_5321_0 = v_5322_0 | v_9301_0;
  assign v_5322_0 = v_5323_0 | v_9300_0;
  assign v_5323_0 = v_589_0 ? v_5324_0 : 3'h0;
  assign v_5325_0 = v_5326_0 | v_5327_0;
  assign v_5326_0 = v_589_0 | v_601_0;
  assign v_5327_0 = v_607_0 | v_26_0;
  assign v_5328_0 = v_5329_0 | v_9297_0;
  assign v_5329_0 = v_5330_0 | v_9296_0;
  assign v_5330_0 = v_589_0 ? v_5331_0 : 3'h0;
  assign v_5332_0 = v_5333_0 | v_5334_0;
  assign v_5333_0 = v_589_0 | v_601_0;
  assign v_5334_0 = v_607_0 | v_26_0;
  assign v_5335_0 = v_5336_0 | v_9293_0;
  assign v_5336_0 = v_5337_0 | v_9292_0;
  assign v_5337_0 = v_589_0 ? v_5338_0 : 3'h0;
  assign v_5339_0 = v_5340_0 | v_5341_0;
  assign v_5340_0 = v_589_0 | v_601_0;
  assign v_5341_0 = v_607_0 | v_26_0;
  assign v_5342_0 = v_5343_0 | v_9289_0;
  assign v_5343_0 = v_5344_0 | v_9288_0;
  assign v_5344_0 = v_589_0 ? v_5345_0 : 3'h0;
  assign v_5346_0 = v_5347_0 | v_5348_0;
  assign v_5347_0 = v_589_0 | v_601_0;
  assign v_5348_0 = v_607_0 | v_26_0;
  assign v_5349_0 = v_5350_0 | v_9285_0;
  assign v_5350_0 = v_5351_0 | v_9284_0;
  assign v_5351_0 = v_589_0 ? v_5352_0 : 3'h0;
  assign v_5353_0 = v_5354_0 | v_5355_0;
  assign v_5354_0 = v_589_0 | v_601_0;
  assign v_5355_0 = v_607_0 | v_26_0;
  assign v_5356_0 = v_5357_0 | v_9281_0;
  assign v_5357_0 = v_5358_0 | v_9280_0;
  assign v_5358_0 = v_589_0 ? v_5359_0 : 3'h0;
  assign v_5360_0 = v_5361_0 | v_5362_0;
  assign v_5361_0 = v_589_0 | v_601_0;
  assign v_5362_0 = v_607_0 | v_26_0;
  assign v_5363_0 = v_5364_0 | v_9277_0;
  assign v_5364_0 = v_5365_0 | v_9276_0;
  assign v_5365_0 = v_589_0 ? v_5366_0 : 3'h0;
  assign v_5367_0 = v_5368_0 | v_5369_0;
  assign v_5368_0 = v_589_0 | v_601_0;
  assign v_5369_0 = v_607_0 | v_26_0;
  assign v_5370_0 = v_5371_0 | v_9273_0;
  assign v_5371_0 = v_5372_0 | v_9272_0;
  assign v_5372_0 = v_589_0 ? v_5373_0 : 3'h0;
  assign v_5374_0 = v_5375_0 | v_5376_0;
  assign v_5375_0 = v_589_0 | v_601_0;
  assign v_5376_0 = v_607_0 | v_26_0;
  assign v_5377_0 = v_5378_0 | v_9269_0;
  assign v_5378_0 = v_5379_0 | v_9268_0;
  assign v_5379_0 = v_589_0 ? v_5380_0 : 3'h0;
  assign v_5381_0 = v_5382_0 | v_5383_0;
  assign v_5382_0 = v_589_0 | v_601_0;
  assign v_5383_0 = v_607_0 | v_26_0;
  assign v_5384_0 = v_5385_0 | v_9265_0;
  assign v_5385_0 = v_5386_0 | v_9264_0;
  assign v_5386_0 = v_589_0 ? v_5387_0 : 3'h0;
  assign v_5388_0 = v_5389_0 | v_5390_0;
  assign v_5389_0 = v_589_0 | v_601_0;
  assign v_5390_0 = v_607_0 | v_26_0;
  assign v_5391_0 = v_5392_0 | v_9261_0;
  assign v_5392_0 = v_5393_0 | v_9260_0;
  assign v_5393_0 = v_589_0 ? v_5394_0 : 3'h0;
  assign v_5395_0 = v_5396_0 | v_5397_0;
  assign v_5396_0 = v_589_0 | v_601_0;
  assign v_5397_0 = v_607_0 | v_26_0;
  assign v_5398_0 = v_5399_0 | v_9257_0;
  assign v_5399_0 = v_5400_0 | v_9256_0;
  assign v_5400_0 = v_589_0 ? v_5401_0 : 3'h0;
  assign v_5402_0 = v_5403_0 | v_5404_0;
  assign v_5403_0 = v_589_0 | v_601_0;
  assign v_5404_0 = v_607_0 | v_26_0;
  assign v_5405_0 = v_5406_0 | v_9253_0;
  assign v_5406_0 = v_5407_0 | v_9252_0;
  assign v_5407_0 = v_589_0 ? v_5408_0 : 3'h0;
  assign v_5409_0 = v_5410_0 | v_5411_0;
  assign v_5410_0 = v_589_0 | v_601_0;
  assign v_5411_0 = v_607_0 | v_26_0;
  assign v_5412_0 = v_5413_0 | v_9249_0;
  assign v_5413_0 = v_5414_0 | v_9248_0;
  assign v_5414_0 = v_589_0 ? v_5415_0 : 3'h0;
  assign v_5416_0 = v_5417_0 | v_5418_0;
  assign v_5417_0 = v_589_0 | v_601_0;
  assign v_5418_0 = v_607_0 | v_26_0;
  assign v_5419_0 = v_5420_0 | v_9245_0;
  assign v_5420_0 = v_5421_0 | v_9244_0;
  assign v_5421_0 = v_589_0 ? v_5422_0 : 3'h0;
  assign v_5423_0 = v_5424_0 | v_5425_0;
  assign v_5424_0 = v_589_0 | v_601_0;
  assign v_5425_0 = v_607_0 | v_26_0;
  assign v_5426_0 = v_5427_0 | v_9241_0;
  assign v_5427_0 = v_5428_0 | v_9240_0;
  assign v_5428_0 = v_589_0 ? v_5429_0 : 3'h0;
  assign v_5430_0 = v_5431_0 | v_5432_0;
  assign v_5431_0 = v_589_0 | v_601_0;
  assign v_5432_0 = v_607_0 | v_26_0;
  assign v_5433_0 = v_5434_0 | v_9237_0;
  assign v_5434_0 = v_5435_0 | v_9236_0;
  assign v_5435_0 = v_589_0 ? v_5436_0 : 3'h0;
  assign v_5437_0 = v_5438_0 | v_5439_0;
  assign v_5438_0 = v_589_0 | v_601_0;
  assign v_5439_0 = v_607_0 | v_26_0;
  assign v_5440_0 = v_5441_0 | v_9233_0;
  assign v_5441_0 = v_5442_0 | v_9232_0;
  assign v_5442_0 = v_589_0 ? v_5443_0 : 3'h0;
  assign v_5444_0 = v_5445_0 | v_5446_0;
  assign v_5445_0 = v_589_0 | v_601_0;
  assign v_5446_0 = v_607_0 | v_26_0;
  assign v_5447_0 = v_5448_0 | v_9229_0;
  assign v_5448_0 = v_5449_0 | v_9228_0;
  assign v_5449_0 = v_589_0 ? v_5450_0 : 3'h0;
  assign v_5451_0 = v_5452_0 | v_5453_0;
  assign v_5452_0 = v_589_0 | v_601_0;
  assign v_5453_0 = v_607_0 | v_26_0;
  assign v_5454_0 = v_5455_0 | v_9225_0;
  assign v_5455_0 = v_5456_0 | v_9224_0;
  assign v_5456_0 = v_589_0 ? v_5457_0 : 3'h0;
  assign v_5458_0 = v_5459_0 | v_5460_0;
  assign v_5459_0 = v_589_0 | v_601_0;
  assign v_5460_0 = v_607_0 | v_26_0;
  assign v_5461_0 = v_5462_0 | v_9221_0;
  assign v_5462_0 = v_5463_0 | v_9220_0;
  assign v_5463_0 = v_589_0 ? v_5464_0 : 3'h0;
  assign v_5465_0 = v_5466_0 | v_5467_0;
  assign v_5466_0 = v_589_0 | v_601_0;
  assign v_5467_0 = v_607_0 | v_26_0;
  assign v_5468_0 = v_5469_0 | v_9217_0;
  assign v_5469_0 = v_5470_0 | v_9216_0;
  assign v_5470_0 = v_589_0 ? v_5471_0 : 3'h0;
  assign v_5472_0 = v_5473_0 | v_5474_0;
  assign v_5473_0 = v_589_0 | v_601_0;
  assign v_5474_0 = v_607_0 | v_26_0;
  assign v_5475_0 = v_5476_0 | v_9213_0;
  assign v_5476_0 = v_5477_0 | v_9212_0;
  assign v_5477_0 = v_589_0 ? v_5478_0 : 3'h0;
  assign v_5479_0 = v_5480_0 | v_5481_0;
  assign v_5480_0 = v_589_0 | v_601_0;
  assign v_5481_0 = v_607_0 | v_26_0;
  assign v_5482_0 = v_5483_0 | v_9209_0;
  assign v_5483_0 = v_5484_0 | v_9208_0;
  assign v_5484_0 = v_589_0 ? v_5485_0 : 3'h0;
  assign v_5486_0 = v_5487_0 | v_5488_0;
  assign v_5487_0 = v_589_0 | v_601_0;
  assign v_5488_0 = v_607_0 | v_26_0;
  assign v_5489_0 = v_5490_0 | v_9205_0;
  assign v_5490_0 = v_5491_0 | v_9204_0;
  assign v_5491_0 = v_589_0 ? v_5492_0 : 3'h0;
  assign v_5493_0 = v_5494_0 | v_5495_0;
  assign v_5494_0 = v_589_0 | v_601_0;
  assign v_5495_0 = v_607_0 | v_26_0;
  assign v_5496_0 = v_5497_0 | v_9201_0;
  assign v_5497_0 = v_5498_0 | v_9200_0;
  assign v_5498_0 = v_589_0 ? v_5499_0 : 3'h0;
  assign v_5500_0 = v_5501_0 | v_5502_0;
  assign v_5501_0 = v_589_0 | v_601_0;
  assign v_5502_0 = v_607_0 | v_26_0;
  assign v_5503_0 = v_5504_0 | v_9197_0;
  assign v_5504_0 = v_5505_0 | v_9196_0;
  assign v_5505_0 = v_589_0 ? v_5506_0 : 3'h0;
  assign v_5507_0 = v_5508_0 | v_5509_0;
  assign v_5508_0 = v_589_0 | v_601_0;
  assign v_5509_0 = v_607_0 | v_26_0;
  assign v_5510_0 = v_5511_0 | v_9193_0;
  assign v_5511_0 = v_5512_0 | v_9192_0;
  assign v_5512_0 = v_589_0 ? v_5513_0 : 3'h0;
  assign v_5514_0 = v_5515_0 | v_5516_0;
  assign v_5515_0 = v_589_0 | v_601_0;
  assign v_5516_0 = v_607_0 | v_26_0;
  assign v_5517_0 = v_5518_0 | v_9189_0;
  assign v_5518_0 = v_5519_0 | v_9188_0;
  assign v_5519_0 = v_589_0 ? v_5520_0 : 3'h0;
  assign v_5521_0 = v_5522_0 | v_5523_0;
  assign v_5522_0 = v_589_0 | v_601_0;
  assign v_5523_0 = v_607_0 | v_26_0;
  assign v_5524_0 = v_5525_0 | v_9185_0;
  assign v_5525_0 = v_5526_0 | v_9184_0;
  assign v_5526_0 = v_589_0 ? v_5527_0 : 3'h0;
  assign v_5528_0 = v_5529_0 | v_5530_0;
  assign v_5529_0 = v_589_0 | v_601_0;
  assign v_5530_0 = v_607_0 | v_26_0;
  assign v_5531_0 = v_5532_0 | v_9181_0;
  assign v_5532_0 = v_5533_0 | v_9180_0;
  assign v_5533_0 = v_589_0 ? v_5534_0 : 3'h0;
  assign v_5535_0 = v_5536_0 | v_5537_0;
  assign v_5536_0 = v_589_0 | v_601_0;
  assign v_5537_0 = v_607_0 | v_26_0;
  assign v_5538_0 = v_5539_0 | v_9177_0;
  assign v_5539_0 = v_5540_0 | v_9176_0;
  assign v_5540_0 = v_589_0 ? v_5541_0 : 3'h0;
  assign v_5542_0 = v_5543_0 | v_5544_0;
  assign v_5543_0 = v_589_0 | v_601_0;
  assign v_5544_0 = v_607_0 | v_26_0;
  assign v_5545_0 = v_5546_0 | v_9173_0;
  assign v_5546_0 = v_5547_0 | v_9172_0;
  assign v_5547_0 = v_589_0 ? v_5548_0 : 3'h0;
  assign v_5549_0 = v_5550_0 | v_5551_0;
  assign v_5550_0 = v_589_0 | v_601_0;
  assign v_5551_0 = v_607_0 | v_26_0;
  assign v_5552_0 = v_5553_0 | v_9169_0;
  assign v_5553_0 = v_5554_0 | v_9168_0;
  assign v_5554_0 = v_589_0 ? v_5555_0 : 3'h0;
  assign v_5556_0 = v_5557_0 | v_5558_0;
  assign v_5557_0 = v_589_0 | v_601_0;
  assign v_5558_0 = v_607_0 | v_26_0;
  assign v_5559_0 = v_5560_0 | v_9165_0;
  assign v_5560_0 = v_5561_0 | v_9164_0;
  assign v_5561_0 = v_589_0 ? v_5562_0 : 3'h0;
  assign v_5563_0 = v_5564_0 | v_5565_0;
  assign v_5564_0 = v_589_0 | v_601_0;
  assign v_5565_0 = v_607_0 | v_26_0;
  assign v_5566_0 = v_5567_0 | v_9161_0;
  assign v_5567_0 = v_5568_0 | v_9160_0;
  assign v_5568_0 = v_589_0 ? v_5569_0 : 3'h0;
  assign v_5570_0 = v_5571_0 | v_5572_0;
  assign v_5571_0 = v_589_0 | v_601_0;
  assign v_5572_0 = v_607_0 | v_26_0;
  assign v_5573_0 = v_5574_0 | v_9157_0;
  assign v_5574_0 = v_5575_0 | v_9156_0;
  assign v_5575_0 = v_589_0 ? v_5576_0 : 3'h0;
  assign v_5577_0 = v_5578_0 | v_5579_0;
  assign v_5578_0 = v_589_0 | v_601_0;
  assign v_5579_0 = v_607_0 | v_26_0;
  assign v_5580_0 = v_5581_0 | v_9153_0;
  assign v_5581_0 = v_5582_0 | v_9152_0;
  assign v_5582_0 = v_589_0 ? v_5583_0 : 3'h0;
  assign v_5584_0 = v_5585_0 | v_5586_0;
  assign v_5585_0 = v_589_0 | v_601_0;
  assign v_5586_0 = v_607_0 | v_26_0;
  assign v_5587_0 = v_5588_0 | v_9149_0;
  assign v_5588_0 = v_5589_0 | v_9148_0;
  assign v_5589_0 = v_589_0 ? v_5590_0 : 3'h0;
  assign v_5591_0 = v_5592_0 | v_5593_0;
  assign v_5592_0 = v_589_0 | v_601_0;
  assign v_5593_0 = v_607_0 | v_26_0;
  assign v_5594_0 = v_5595_0 | v_9145_0;
  assign v_5595_0 = v_5596_0 | v_9144_0;
  assign v_5596_0 = v_589_0 ? v_5597_0 : 3'h0;
  assign v_5598_0 = v_5599_0 | v_5600_0;
  assign v_5599_0 = v_589_0 | v_601_0;
  assign v_5600_0 = v_607_0 | v_26_0;
  assign v_5601_0 = v_5602_0 | v_9141_0;
  assign v_5602_0 = v_5603_0 | v_9140_0;
  assign v_5603_0 = v_589_0 ? v_5604_0 : 3'h0;
  assign v_5605_0 = v_5606_0 | v_5607_0;
  assign v_5606_0 = v_589_0 | v_601_0;
  assign v_5607_0 = v_607_0 | v_26_0;
  assign v_5608_0 = v_5609_0 | v_9137_0;
  assign v_5609_0 = v_5610_0 | v_9136_0;
  assign v_5610_0 = v_589_0 ? v_5611_0 : 3'h0;
  assign v_5612_0 = v_5613_0 | v_5614_0;
  assign v_5613_0 = v_589_0 | v_601_0;
  assign v_5614_0 = v_607_0 | v_26_0;
  assign v_5615_0 = v_5616_0 | v_9133_0;
  assign v_5616_0 = v_5617_0 | v_9132_0;
  assign v_5617_0 = v_589_0 ? v_5618_0 : 3'h0;
  assign v_5619_0 = v_5620_0 | v_5621_0;
  assign v_5620_0 = v_589_0 | v_601_0;
  assign v_5621_0 = v_607_0 | v_26_0;
  assign v_5622_0 = v_5623_0 | v_9129_0;
  assign v_5623_0 = v_5624_0 | v_9128_0;
  assign v_5624_0 = v_589_0 ? v_5625_0 : 3'h0;
  assign v_5626_0 = v_5627_0 | v_5628_0;
  assign v_5627_0 = v_589_0 | v_601_0;
  assign v_5628_0 = v_607_0 | v_26_0;
  assign v_5629_0 = v_5630_0 | v_9125_0;
  assign v_5630_0 = v_5631_0 | v_9124_0;
  assign v_5631_0 = v_589_0 ? v_5632_0 : 3'h0;
  assign v_5633_0 = v_5634_0 | v_5635_0;
  assign v_5634_0 = v_589_0 | v_601_0;
  assign v_5635_0 = v_607_0 | v_26_0;
  assign v_5636_0 = v_5637_0 | v_9121_0;
  assign v_5637_0 = v_5638_0 | v_9120_0;
  assign v_5638_0 = v_589_0 ? v_5639_0 : 3'h0;
  assign v_5640_0 = v_5641_0 | v_5642_0;
  assign v_5641_0 = v_589_0 | v_601_0;
  assign v_5642_0 = v_607_0 | v_26_0;
  assign v_5643_0 = v_5644_0 | v_9117_0;
  assign v_5644_0 = v_5645_0 | v_9116_0;
  assign v_5645_0 = v_589_0 ? v_5646_0 : 3'h0;
  assign v_5647_0 = v_5648_0 | v_5649_0;
  assign v_5648_0 = v_589_0 | v_601_0;
  assign v_5649_0 = v_607_0 | v_26_0;
  assign v_5650_0 = v_5651_0 | v_9113_0;
  assign v_5651_0 = v_5652_0 | v_9112_0;
  assign v_5652_0 = v_589_0 ? v_5653_0 : 3'h0;
  assign v_5654_0 = v_5655_0 | v_5656_0;
  assign v_5655_0 = v_589_0 | v_601_0;
  assign v_5656_0 = v_607_0 | v_26_0;
  assign v_5657_0 = v_5658_0 | v_9109_0;
  assign v_5658_0 = v_5659_0 | v_9108_0;
  assign v_5659_0 = v_589_0 ? v_5660_0 : 3'h0;
  assign v_5661_0 = v_5662_0 | v_5663_0;
  assign v_5662_0 = v_589_0 | v_601_0;
  assign v_5663_0 = v_607_0 | v_26_0;
  assign v_5664_0 = v_5665_0 | v_9105_0;
  assign v_5665_0 = v_5666_0 | v_9104_0;
  assign v_5666_0 = v_589_0 ? v_5667_0 : 3'h0;
  assign v_5668_0 = v_5669_0 | v_5670_0;
  assign v_5669_0 = v_589_0 | v_601_0;
  assign v_5670_0 = v_607_0 | v_26_0;
  assign v_5671_0 = v_5672_0 | v_9101_0;
  assign v_5672_0 = v_5673_0 | v_9100_0;
  assign v_5673_0 = v_589_0 ? v_5674_0 : 3'h0;
  assign v_5675_0 = v_5676_0 | v_5677_0;
  assign v_5676_0 = v_589_0 | v_601_0;
  assign v_5677_0 = v_607_0 | v_26_0;
  assign v_5678_0 = v_5679_0 | v_9097_0;
  assign v_5679_0 = v_5680_0 | v_9096_0;
  assign v_5680_0 = v_589_0 ? v_5681_0 : 3'h0;
  assign v_5682_0 = v_5683_0 | v_5684_0;
  assign v_5683_0 = v_589_0 | v_601_0;
  assign v_5684_0 = v_607_0 | v_26_0;
  assign v_5685_0 = v_5686_0 | v_9093_0;
  assign v_5686_0 = v_5687_0 | v_9092_0;
  assign v_5687_0 = v_589_0 ? v_5688_0 : 3'h0;
  assign v_5689_0 = v_5690_0 | v_5691_0;
  assign v_5690_0 = v_589_0 | v_601_0;
  assign v_5691_0 = v_607_0 | v_26_0;
  assign v_5692_0 = v_5693_0 | v_9089_0;
  assign v_5693_0 = v_5694_0 | v_9088_0;
  assign v_5694_0 = v_589_0 ? v_5695_0 : 3'h0;
  assign v_5696_0 = v_5697_0 | v_5698_0;
  assign v_5697_0 = v_589_0 | v_601_0;
  assign v_5698_0 = v_607_0 | v_26_0;
  assign v_5699_0 = v_5700_0 | v_9085_0;
  assign v_5700_0 = v_5701_0 | v_9084_0;
  assign v_5701_0 = v_589_0 ? v_5702_0 : 3'h0;
  assign v_5703_0 = v_5704_0 | v_5705_0;
  assign v_5704_0 = v_589_0 | v_601_0;
  assign v_5705_0 = v_607_0 | v_26_0;
  assign v_5706_0 = v_5707_0 | v_9081_0;
  assign v_5707_0 = v_5708_0 | v_9080_0;
  assign v_5708_0 = v_589_0 ? v_5709_0 : 3'h0;
  assign v_5710_0 = v_5711_0 | v_5712_0;
  assign v_5711_0 = v_589_0 | v_601_0;
  assign v_5712_0 = v_607_0 | v_26_0;
  assign v_5713_0 = v_5714_0 | v_9077_0;
  assign v_5714_0 = v_5715_0 | v_9076_0;
  assign v_5715_0 = v_589_0 ? v_5716_0 : 3'h0;
  assign v_5717_0 = v_5718_0 | v_5719_0;
  assign v_5718_0 = v_589_0 | v_601_0;
  assign v_5719_0 = v_607_0 | v_26_0;
  assign v_5720_0 = v_5721_0 | v_9073_0;
  assign v_5721_0 = v_5722_0 | v_9072_0;
  assign v_5722_0 = v_589_0 ? v_5723_0 : 3'h0;
  assign v_5724_0 = v_5725_0 | v_5726_0;
  assign v_5725_0 = v_589_0 | v_601_0;
  assign v_5726_0 = v_607_0 | v_26_0;
  assign v_5727_0 = v_5728_0 | v_9069_0;
  assign v_5728_0 = v_5729_0 | v_9068_0;
  assign v_5729_0 = v_589_0 ? v_5730_0 : 3'h0;
  assign v_5731_0 = v_5732_0 | v_5733_0;
  assign v_5732_0 = v_589_0 | v_601_0;
  assign v_5733_0 = v_607_0 | v_26_0;
  assign v_5734_0 = v_5735_0 | v_9065_0;
  assign v_5735_0 = v_5736_0 | v_9064_0;
  assign v_5736_0 = v_589_0 ? v_5737_0 : 3'h0;
  assign v_5738_0 = v_5739_0 | v_5740_0;
  assign v_5739_0 = v_589_0 | v_601_0;
  assign v_5740_0 = v_607_0 | v_26_0;
  assign v_5741_0 = v_5742_0 | v_9061_0;
  assign v_5742_0 = v_5743_0 | v_9060_0;
  assign v_5743_0 = v_589_0 ? v_5744_0 : 3'h0;
  assign v_5745_0 = v_5746_0 | v_5747_0;
  assign v_5746_0 = v_589_0 | v_601_0;
  assign v_5747_0 = v_607_0 | v_26_0;
  assign v_5748_0 = v_5749_0 | v_9057_0;
  assign v_5749_0 = v_5750_0 | v_9056_0;
  assign v_5750_0 = v_589_0 ? v_5751_0 : 3'h0;
  assign v_5752_0 = v_5753_0 | v_5754_0;
  assign v_5753_0 = v_589_0 | v_601_0;
  assign v_5754_0 = v_607_0 | v_26_0;
  assign v_5755_0 = v_5756_0 | v_9053_0;
  assign v_5756_0 = v_5757_0 | v_9052_0;
  assign v_5757_0 = v_589_0 ? v_5758_0 : 3'h0;
  assign v_5759_0 = v_5760_0 | v_5761_0;
  assign v_5760_0 = v_589_0 | v_601_0;
  assign v_5761_0 = v_607_0 | v_26_0;
  assign v_5762_0 = v_5763_0 | v_9049_0;
  assign v_5763_0 = v_5764_0 | v_9048_0;
  assign v_5764_0 = v_589_0 ? v_5765_0 : 3'h0;
  assign v_5766_0 = v_5767_0 | v_5768_0;
  assign v_5767_0 = v_589_0 | v_601_0;
  assign v_5768_0 = v_607_0 | v_26_0;
  assign v_5769_0 = v_5770_0 | v_9045_0;
  assign v_5770_0 = v_5771_0 | v_9044_0;
  assign v_5771_0 = v_589_0 ? v_5772_0 : 3'h0;
  assign v_5773_0 = v_5774_0 | v_5775_0;
  assign v_5774_0 = v_589_0 | v_601_0;
  assign v_5775_0 = v_607_0 | v_26_0;
  assign v_5776_0 = v_5777_0 | v_9041_0;
  assign v_5777_0 = v_5778_0 | v_9040_0;
  assign v_5778_0 = v_589_0 ? v_5779_0 : 3'h0;
  assign v_5780_0 = v_5781_0 | v_5782_0;
  assign v_5781_0 = v_589_0 | v_601_0;
  assign v_5782_0 = v_607_0 | v_26_0;
  assign v_5783_0 = v_5784_0 | v_9037_0;
  assign v_5784_0 = v_5785_0 | v_9036_0;
  assign v_5785_0 = v_589_0 ? v_5786_0 : 3'h0;
  assign v_5787_0 = v_5788_0 | v_5789_0;
  assign v_5788_0 = v_589_0 | v_601_0;
  assign v_5789_0 = v_607_0 | v_26_0;
  assign v_5790_0 = v_5791_0 | v_9033_0;
  assign v_5791_0 = v_5792_0 | v_9032_0;
  assign v_5792_0 = v_589_0 ? v_5793_0 : 3'h0;
  assign v_5794_0 = v_5795_0 | v_5796_0;
  assign v_5795_0 = v_589_0 | v_601_0;
  assign v_5796_0 = v_607_0 | v_26_0;
  assign v_5797_0 = v_5798_0 | v_9029_0;
  assign v_5798_0 = v_5799_0 | v_9028_0;
  assign v_5799_0 = v_589_0 ? v_5800_0 : 3'h0;
  assign v_5801_0 = v_5802_0 | v_5803_0;
  assign v_5802_0 = v_589_0 | v_601_0;
  assign v_5803_0 = v_607_0 | v_26_0;
  assign v_5804_0 = v_5805_0 | v_9025_0;
  assign v_5805_0 = v_5806_0 | v_9024_0;
  assign v_5806_0 = v_589_0 ? v_5807_0 : 3'h0;
  assign v_5808_0 = v_5809_0 | v_5810_0;
  assign v_5809_0 = v_589_0 | v_601_0;
  assign v_5810_0 = v_607_0 | v_26_0;
  assign v_5811_0 = v_5812_0 | v_9021_0;
  assign v_5812_0 = v_5813_0 | v_9020_0;
  assign v_5813_0 = v_589_0 ? v_5814_0 : 3'h0;
  assign v_5815_0 = v_5816_0 | v_5817_0;
  assign v_5816_0 = v_589_0 | v_601_0;
  assign v_5817_0 = v_607_0 | v_26_0;
  assign v_5818_0 = v_5819_0 | v_9017_0;
  assign v_5819_0 = v_5820_0 | v_9016_0;
  assign v_5820_0 = v_589_0 ? v_5821_0 : 3'h0;
  assign v_5822_0 = v_5823_0 | v_5824_0;
  assign v_5823_0 = v_589_0 | v_601_0;
  assign v_5824_0 = v_607_0 | v_26_0;
  assign v_5825_0 = v_5826_0 | v_9013_0;
  assign v_5826_0 = v_5827_0 | v_9012_0;
  assign v_5827_0 = v_589_0 ? v_5828_0 : 3'h0;
  assign v_5829_0 = v_5830_0 | v_5831_0;
  assign v_5830_0 = v_589_0 | v_601_0;
  assign v_5831_0 = v_607_0 | v_26_0;
  assign v_5832_0 = v_5833_0 | v_9009_0;
  assign v_5833_0 = v_5834_0 | v_9008_0;
  assign v_5834_0 = v_589_0 ? v_5835_0 : 3'h0;
  assign v_5836_0 = v_5837_0 | v_5838_0;
  assign v_5837_0 = v_589_0 | v_601_0;
  assign v_5838_0 = v_607_0 | v_26_0;
  assign v_5839_0 = v_5840_0 | v_9005_0;
  assign v_5840_0 = v_5841_0 | v_9004_0;
  assign v_5841_0 = v_589_0 ? v_5842_0 : 3'h0;
  assign v_5843_0 = v_5844_0 | v_5845_0;
  assign v_5844_0 = v_589_0 | v_601_0;
  assign v_5845_0 = v_607_0 | v_26_0;
  assign v_5846_0 = v_5847_0 | v_9001_0;
  assign v_5847_0 = v_5848_0 | v_9000_0;
  assign v_5848_0 = v_589_0 ? v_5849_0 : 3'h0;
  assign v_5850_0 = v_5851_0 | v_5852_0;
  assign v_5851_0 = v_589_0 | v_601_0;
  assign v_5852_0 = v_607_0 | v_26_0;
  assign v_5853_0 = v_5854_0 | v_8997_0;
  assign v_5854_0 = v_5855_0 | v_8996_0;
  assign v_5855_0 = v_589_0 ? v_5856_0 : 3'h0;
  assign v_5857_0 = v_5858_0 | v_5859_0;
  assign v_5858_0 = v_589_0 | v_601_0;
  assign v_5859_0 = v_607_0 | v_26_0;
  assign v_5860_0 = v_5861_0 | v_8993_0;
  assign v_5861_0 = v_5862_0 | v_8992_0;
  assign v_5862_0 = v_589_0 ? v_5863_0 : 3'h0;
  assign v_5864_0 = v_5865_0 | v_5866_0;
  assign v_5865_0 = v_589_0 | v_601_0;
  assign v_5866_0 = v_607_0 | v_26_0;
  assign v_5867_0 = v_5868_0 | v_8989_0;
  assign v_5868_0 = v_5869_0 | v_8988_0;
  assign v_5869_0 = v_589_0 ? v_5870_0 : 3'h0;
  assign v_5871_0 = v_5872_0 | v_5873_0;
  assign v_5872_0 = v_589_0 | v_601_0;
  assign v_5873_0 = v_607_0 | v_26_0;
  assign v_5874_0 = v_5875_0 | v_8985_0;
  assign v_5875_0 = v_5876_0 | v_8984_0;
  assign v_5876_0 = v_589_0 ? v_5877_0 : 3'h0;
  assign v_5878_0 = v_5879_0 | v_5880_0;
  assign v_5879_0 = v_589_0 | v_601_0;
  assign v_5880_0 = v_607_0 | v_26_0;
  assign v_5881_0 = v_5882_0 | v_8981_0;
  assign v_5882_0 = v_5883_0 | v_8980_0;
  assign v_5883_0 = v_589_0 ? v_5884_0 : 3'h0;
  assign v_5885_0 = v_5886_0 | v_5887_0;
  assign v_5886_0 = v_589_0 | v_601_0;
  assign v_5887_0 = v_607_0 | v_26_0;
  assign v_5888_0 = v_5889_0 | v_8977_0;
  assign v_5889_0 = v_5890_0 | v_8976_0;
  assign v_5890_0 = v_589_0 ? v_5891_0 : 3'h0;
  assign v_5892_0 = v_5893_0 | v_5894_0;
  assign v_5893_0 = v_589_0 | v_601_0;
  assign v_5894_0 = v_607_0 | v_26_0;
  assign v_5895_0 = v_5896_0 | v_8973_0;
  assign v_5896_0 = v_5897_0 | v_8972_0;
  assign v_5897_0 = v_589_0 ? v_5898_0 : 3'h0;
  assign v_5899_0 = v_5900_0 | v_5901_0;
  assign v_5900_0 = v_589_0 | v_601_0;
  assign v_5901_0 = v_607_0 | v_26_0;
  assign v_5902_0 = v_5903_0 | v_8969_0;
  assign v_5903_0 = v_5904_0 | v_8968_0;
  assign v_5904_0 = v_589_0 ? v_5905_0 : 3'h0;
  assign v_5906_0 = v_5907_0 | v_5908_0;
  assign v_5907_0 = v_589_0 | v_601_0;
  assign v_5908_0 = v_607_0 | v_26_0;
  assign v_5909_0 = v_5910_0 | v_8965_0;
  assign v_5910_0 = v_5911_0 | v_8964_0;
  assign v_5911_0 = v_589_0 ? v_5912_0 : 3'h0;
  assign v_5913_0 = v_5914_0 | v_5915_0;
  assign v_5914_0 = v_589_0 | v_601_0;
  assign v_5915_0 = v_607_0 | v_26_0;
  assign v_5916_0 = v_5917_0 | v_8961_0;
  assign v_5917_0 = v_5918_0 | v_8960_0;
  assign v_5918_0 = v_589_0 ? v_5919_0 : 3'h0;
  assign v_5920_0 = v_5921_0 | v_5922_0;
  assign v_5921_0 = v_589_0 | v_601_0;
  assign v_5922_0 = v_607_0 | v_26_0;
  assign v_5923_0 = v_5924_0 | v_8957_0;
  assign v_5924_0 = v_5925_0 | v_8956_0;
  assign v_5925_0 = v_589_0 ? v_5926_0 : 3'h0;
  assign v_5927_0 = v_5928_0 | v_5929_0;
  assign v_5928_0 = v_589_0 | v_601_0;
  assign v_5929_0 = v_607_0 | v_26_0;
  assign v_5930_0 = v_5931_0 | v_8953_0;
  assign v_5931_0 = v_5932_0 | v_8952_0;
  assign v_5932_0 = v_589_0 ? v_5933_0 : 3'h0;
  assign v_5934_0 = v_5935_0 | v_5936_0;
  assign v_5935_0 = v_589_0 | v_601_0;
  assign v_5936_0 = v_607_0 | v_26_0;
  assign v_5937_0 = v_5938_0 | v_8949_0;
  assign v_5938_0 = v_5939_0 | v_8948_0;
  assign v_5939_0 = v_589_0 ? v_5940_0 : 3'h0;
  assign v_5941_0 = v_5942_0 | v_5943_0;
  assign v_5942_0 = v_589_0 | v_601_0;
  assign v_5943_0 = v_607_0 | v_26_0;
  assign v_5944_0 = v_5945_0 | v_8945_0;
  assign v_5945_0 = v_5946_0 | v_8944_0;
  assign v_5946_0 = v_589_0 ? v_5947_0 : 3'h0;
  assign v_5948_0 = v_5949_0 | v_5950_0;
  assign v_5949_0 = v_589_0 | v_601_0;
  assign v_5950_0 = v_607_0 | v_26_0;
  assign v_5951_0 = v_5952_0 | v_8941_0;
  assign v_5952_0 = v_5953_0 | v_8940_0;
  assign v_5953_0 = v_589_0 ? v_5954_0 : 3'h0;
  assign v_5955_0 = v_5956_0 | v_5957_0;
  assign v_5956_0 = v_589_0 | v_601_0;
  assign v_5957_0 = v_607_0 | v_26_0;
  assign v_5958_0 = v_5959_0 | v_8937_0;
  assign v_5959_0 = v_5960_0 | v_8936_0;
  assign v_5960_0 = v_589_0 ? v_5961_0 : 3'h0;
  assign v_5962_0 = v_5963_0 | v_5964_0;
  assign v_5963_0 = v_589_0 | v_601_0;
  assign v_5964_0 = v_607_0 | v_26_0;
  assign v_5965_0 = v_5966_0 | v_8933_0;
  assign v_5966_0 = v_5967_0 | v_8932_0;
  assign v_5967_0 = v_589_0 ? v_5968_0 : 3'h0;
  assign v_5969_0 = v_5970_0 | v_5971_0;
  assign v_5970_0 = v_589_0 | v_601_0;
  assign v_5971_0 = v_607_0 | v_26_0;
  assign v_5972_0 = v_5973_0 | v_8929_0;
  assign v_5973_0 = v_5974_0 | v_8928_0;
  assign v_5974_0 = v_589_0 ? v_5975_0 : 3'h0;
  assign v_5976_0 = v_5977_0 | v_5978_0;
  assign v_5977_0 = v_589_0 | v_601_0;
  assign v_5978_0 = v_607_0 | v_26_0;
  assign v_5979_0 = v_5980_0 | v_8925_0;
  assign v_5980_0 = v_5981_0 | v_8924_0;
  assign v_5981_0 = v_589_0 ? v_5982_0 : 3'h0;
  assign v_5983_0 = v_5984_0 | v_5985_0;
  assign v_5984_0 = v_589_0 | v_601_0;
  assign v_5985_0 = v_607_0 | v_26_0;
  assign v_5986_0 = v_5987_0 | v_8921_0;
  assign v_5987_0 = v_5988_0 | v_8920_0;
  assign v_5988_0 = v_589_0 ? v_5989_0 : 3'h0;
  assign v_5990_0 = v_5991_0 | v_5992_0;
  assign v_5991_0 = v_589_0 | v_601_0;
  assign v_5992_0 = v_607_0 | v_26_0;
  assign v_5993_0 = v_5994_0 | v_8917_0;
  assign v_5994_0 = v_5995_0 | v_8916_0;
  assign v_5995_0 = v_589_0 ? v_5996_0 : 3'h0;
  assign v_5997_0 = v_5998_0 | v_5999_0;
  assign v_5998_0 = v_589_0 | v_601_0;
  assign v_5999_0 = v_607_0 | v_26_0;
  assign v_6000_0 = v_6001_0 | v_8913_0;
  assign v_6001_0 = v_6002_0 | v_8912_0;
  assign v_6002_0 = v_589_0 ? v_6003_0 : 3'h0;
  assign v_6004_0 = v_6005_0 | v_6006_0;
  assign v_6005_0 = v_589_0 | v_601_0;
  assign v_6006_0 = v_607_0 | v_26_0;
  assign v_6007_0 = v_6008_0 | v_8909_0;
  assign v_6008_0 = v_6009_0 | v_8908_0;
  assign v_6009_0 = v_589_0 ? v_6010_0 : 3'h0;
  assign v_6011_0 = v_6012_0 | v_6013_0;
  assign v_6012_0 = v_589_0 | v_601_0;
  assign v_6013_0 = v_607_0 | v_26_0;
  assign v_6014_0 = v_6015_0 | v_8905_0;
  assign v_6015_0 = v_6016_0 | v_8904_0;
  assign v_6016_0 = v_589_0 ? v_6017_0 : 3'h0;
  assign v_6018_0 = v_6019_0 | v_6020_0;
  assign v_6019_0 = v_589_0 | v_601_0;
  assign v_6020_0 = v_607_0 | v_26_0;
  assign v_6021_0 = v_6022_0 | v_8901_0;
  assign v_6022_0 = v_6023_0 | v_8900_0;
  assign v_6023_0 = v_589_0 ? v_6024_0 : 3'h0;
  assign v_6025_0 = v_6026_0 | v_6027_0;
  assign v_6026_0 = v_589_0 | v_601_0;
  assign v_6027_0 = v_607_0 | v_26_0;
  assign v_6028_0 = v_6029_0 | v_8897_0;
  assign v_6029_0 = v_6030_0 | v_8896_0;
  assign v_6030_0 = v_589_0 ? v_6031_0 : 3'h0;
  assign v_6032_0 = v_6033_0 | v_6034_0;
  assign v_6033_0 = v_589_0 | v_601_0;
  assign v_6034_0 = v_607_0 | v_26_0;
  assign v_6035_0 = v_6036_0 | v_8893_0;
  assign v_6036_0 = v_6037_0 | v_8892_0;
  assign v_6037_0 = v_589_0 ? v_6038_0 : 3'h0;
  assign v_6039_0 = v_6040_0 | v_6041_0;
  assign v_6040_0 = v_589_0 | v_601_0;
  assign v_6041_0 = v_607_0 | v_26_0;
  assign v_6042_0 = v_6043_0 | v_8889_0;
  assign v_6043_0 = v_6044_0 | v_8888_0;
  assign v_6044_0 = v_589_0 ? v_6045_0 : 3'h0;
  assign v_6046_0 = v_6047_0 | v_6048_0;
  assign v_6047_0 = v_589_0 | v_601_0;
  assign v_6048_0 = v_607_0 | v_26_0;
  assign v_6049_0 = v_6050_0 | v_8885_0;
  assign v_6050_0 = v_6051_0 | v_8884_0;
  assign v_6051_0 = v_589_0 ? v_6052_0 : 3'h0;
  assign v_6053_0 = v_6054_0 | v_6055_0;
  assign v_6054_0 = v_589_0 | v_601_0;
  assign v_6055_0 = v_607_0 | v_26_0;
  assign v_6056_0 = v_6057_0 | v_8881_0;
  assign v_6057_0 = v_6058_0 | v_8880_0;
  assign v_6058_0 = v_589_0 ? v_6059_0 : 3'h0;
  assign v_6060_0 = v_6061_0 | v_6062_0;
  assign v_6061_0 = v_589_0 | v_601_0;
  assign v_6062_0 = v_607_0 | v_26_0;
  assign v_6063_0 = v_6064_0 | v_8877_0;
  assign v_6064_0 = v_6065_0 | v_8876_0;
  assign v_6065_0 = v_589_0 ? v_6066_0 : 3'h0;
  assign v_6067_0 = v_6068_0 | v_6069_0;
  assign v_6068_0 = v_589_0 | v_601_0;
  assign v_6069_0 = v_607_0 | v_26_0;
  assign v_6070_0 = v_6071_0 | v_8873_0;
  assign v_6071_0 = v_6072_0 | v_8872_0;
  assign v_6072_0 = v_589_0 ? v_6073_0 : 3'h0;
  assign v_6074_0 = v_6075_0 | v_6076_0;
  assign v_6075_0 = v_589_0 | v_601_0;
  assign v_6076_0 = v_607_0 | v_26_0;
  assign v_6077_0 = v_6078_0 | v_8869_0;
  assign v_6078_0 = v_6079_0 | v_8868_0;
  assign v_6079_0 = v_589_0 ? v_6080_0 : 3'h0;
  assign v_6081_0 = v_6082_0 | v_6083_0;
  assign v_6082_0 = v_589_0 | v_601_0;
  assign v_6083_0 = v_607_0 | v_26_0;
  assign v_6084_0 = v_6085_0 | v_8865_0;
  assign v_6085_0 = v_6086_0 | v_8864_0;
  assign v_6086_0 = v_589_0 ? v_6087_0 : 3'h0;
  assign v_6088_0 = v_6089_0 | v_6090_0;
  assign v_6089_0 = v_589_0 | v_601_0;
  assign v_6090_0 = v_607_0 | v_26_0;
  assign v_6091_0 = v_6092_0 | v_8861_0;
  assign v_6092_0 = v_6093_0 | v_8860_0;
  assign v_6093_0 = v_589_0 ? v_6094_0 : 3'h0;
  assign v_6095_0 = v_6096_0 | v_6097_0;
  assign v_6096_0 = v_589_0 | v_601_0;
  assign v_6097_0 = v_607_0 | v_26_0;
  assign v_6098_0 = v_6099_0 | v_8857_0;
  assign v_6099_0 = v_6100_0 | v_8856_0;
  assign v_6100_0 = v_589_0 ? v_6101_0 : 3'h0;
  assign v_6102_0 = v_6103_0 | v_6104_0;
  assign v_6103_0 = v_589_0 | v_601_0;
  assign v_6104_0 = v_607_0 | v_26_0;
  assign v_6105_0 = v_6106_0 | v_8853_0;
  assign v_6106_0 = v_6107_0 | v_8852_0;
  assign v_6107_0 = v_589_0 ? v_6108_0 : 3'h0;
  assign v_6109_0 = v_6110_0 | v_6111_0;
  assign v_6110_0 = v_589_0 | v_601_0;
  assign v_6111_0 = v_607_0 | v_26_0;
  assign v_6112_0 = v_6113_0 | v_8849_0;
  assign v_6113_0 = v_6114_0 | v_8848_0;
  assign v_6114_0 = v_589_0 ? v_6115_0 : 3'h0;
  assign v_6116_0 = v_6117_0 | v_6118_0;
  assign v_6117_0 = v_589_0 | v_601_0;
  assign v_6118_0 = v_607_0 | v_26_0;
  assign v_6119_0 = v_6120_0 | v_8845_0;
  assign v_6120_0 = v_6121_0 | v_8844_0;
  assign v_6121_0 = v_589_0 ? v_6122_0 : 3'h0;
  assign v_6123_0 = v_6124_0 | v_6125_0;
  assign v_6124_0 = v_589_0 | v_601_0;
  assign v_6125_0 = v_607_0 | v_26_0;
  assign v_6126_0 = v_6127_0 | v_8841_0;
  assign v_6127_0 = v_6128_0 | v_8840_0;
  assign v_6128_0 = v_589_0 ? v_6129_0 : 3'h0;
  assign v_6130_0 = v_6131_0 | v_6132_0;
  assign v_6131_0 = v_589_0 | v_601_0;
  assign v_6132_0 = v_607_0 | v_26_0;
  assign v_6133_0 = v_6134_0 | v_8837_0;
  assign v_6134_0 = v_6135_0 | v_8836_0;
  assign v_6135_0 = v_589_0 ? v_6136_0 : 3'h0;
  assign v_6137_0 = v_6138_0 | v_6139_0;
  assign v_6138_0 = v_589_0 | v_601_0;
  assign v_6139_0 = v_607_0 | v_26_0;
  assign v_6140_0 = v_6141_0 | v_8833_0;
  assign v_6141_0 = v_6142_0 | v_8832_0;
  assign v_6142_0 = v_589_0 ? v_6143_0 : 3'h0;
  assign v_6144_0 = v_6145_0 | v_6146_0;
  assign v_6145_0 = v_589_0 | v_601_0;
  assign v_6146_0 = v_607_0 | v_26_0;
  assign v_6147_0 = v_6148_0 | v_8829_0;
  assign v_6148_0 = v_6149_0 | v_8828_0;
  assign v_6149_0 = v_589_0 ? v_6150_0 : 3'h0;
  assign v_6151_0 = v_6152_0 | v_6153_0;
  assign v_6152_0 = v_589_0 | v_601_0;
  assign v_6153_0 = v_607_0 | v_26_0;
  assign v_6154_0 = v_6155_0 | v_8825_0;
  assign v_6155_0 = v_6156_0 | v_8824_0;
  assign v_6156_0 = v_589_0 ? v_6157_0 : 3'h0;
  assign v_6158_0 = v_6159_0 | v_6160_0;
  assign v_6159_0 = v_589_0 | v_601_0;
  assign v_6160_0 = v_607_0 | v_26_0;
  assign v_6161_0 = v_6162_0 | v_8821_0;
  assign v_6162_0 = v_6163_0 | v_8820_0;
  assign v_6163_0 = v_589_0 ? v_6164_0 : 3'h0;
  assign v_6165_0 = v_6166_0 | v_6167_0;
  assign v_6166_0 = v_589_0 | v_601_0;
  assign v_6167_0 = v_607_0 | v_26_0;
  assign v_6168_0 = v_6169_0 | v_8817_0;
  assign v_6169_0 = v_6170_0 | v_8816_0;
  assign v_6170_0 = v_589_0 ? v_6171_0 : 3'h0;
  assign v_6172_0 = v_6173_0 | v_6174_0;
  assign v_6173_0 = v_589_0 | v_601_0;
  assign v_6174_0 = v_607_0 | v_26_0;
  assign v_6175_0 = v_6176_0 | v_8813_0;
  assign v_6176_0 = v_6177_0 | v_8812_0;
  assign v_6177_0 = v_589_0 ? v_6178_0 : 3'h0;
  assign v_6179_0 = v_6180_0 | v_6181_0;
  assign v_6180_0 = v_589_0 | v_601_0;
  assign v_6181_0 = v_607_0 | v_26_0;
  assign v_6182_0 = v_6183_0 | v_8809_0;
  assign v_6183_0 = v_6184_0 | v_8808_0;
  assign v_6184_0 = v_589_0 ? v_6185_0 : 3'h0;
  assign v_6186_0 = v_6187_0 | v_6188_0;
  assign v_6187_0 = v_589_0 | v_601_0;
  assign v_6188_0 = v_607_0 | v_26_0;
  assign v_6189_0 = v_6190_0 | v_8805_0;
  assign v_6190_0 = v_6191_0 | v_8804_0;
  assign v_6191_0 = v_589_0 ? v_6192_0 : 3'h0;
  assign v_6193_0 = v_6194_0 | v_6195_0;
  assign v_6194_0 = v_589_0 | v_601_0;
  assign v_6195_0 = v_607_0 | v_26_0;
  assign v_6196_0 = v_6197_0 | v_8801_0;
  assign v_6197_0 = v_6198_0 | v_8800_0;
  assign v_6198_0 = v_589_0 ? v_6199_0 : 3'h0;
  assign v_6200_0 = v_6201_0 | v_6202_0;
  assign v_6201_0 = v_589_0 | v_601_0;
  assign v_6202_0 = v_607_0 | v_26_0;
  assign v_6203_0 = v_6204_0 | v_8797_0;
  assign v_6204_0 = v_6205_0 | v_8796_0;
  assign v_6205_0 = v_589_0 ? v_6206_0 : 3'h0;
  assign v_6207_0 = v_6208_0 | v_6209_0;
  assign v_6208_0 = v_589_0 | v_601_0;
  assign v_6209_0 = v_607_0 | v_26_0;
  assign v_6210_0 = v_6211_0 | v_8793_0;
  assign v_6211_0 = v_6212_0 | v_8792_0;
  assign v_6212_0 = v_589_0 ? v_6213_0 : 3'h0;
  assign v_6214_0 = v_6215_0 | v_6216_0;
  assign v_6215_0 = v_589_0 | v_601_0;
  assign v_6216_0 = v_607_0 | v_26_0;
  assign v_6217_0 = v_6218_0 | v_8789_0;
  assign v_6218_0 = v_6219_0 | v_8788_0;
  assign v_6219_0 = v_589_0 ? v_6220_0 : 3'h0;
  assign v_6221_0 = v_6222_0 | v_6223_0;
  assign v_6222_0 = v_589_0 | v_601_0;
  assign v_6223_0 = v_607_0 | v_26_0;
  assign v_6224_0 = v_6225_0 | v_8785_0;
  assign v_6225_0 = v_6226_0 | v_8784_0;
  assign v_6226_0 = v_589_0 ? v_6227_0 : 3'h0;
  assign v_6228_0 = v_6229_0 | v_6230_0;
  assign v_6229_0 = v_589_0 | v_601_0;
  assign v_6230_0 = v_607_0 | v_26_0;
  assign v_6231_0 = v_6232_0 | v_8781_0;
  assign v_6232_0 = v_6233_0 | v_8780_0;
  assign v_6233_0 = v_589_0 ? v_6234_0 : 3'h0;
  assign v_6235_0 = v_6236_0 | v_6237_0;
  assign v_6236_0 = v_589_0 | v_601_0;
  assign v_6237_0 = v_607_0 | v_26_0;
  assign v_6238_0 = v_6239_0 | v_8777_0;
  assign v_6239_0 = v_6240_0 | v_8776_0;
  assign v_6240_0 = v_589_0 ? v_6241_0 : 3'h0;
  assign v_6242_0 = v_6243_0 | v_6244_0;
  assign v_6243_0 = v_589_0 | v_601_0;
  assign v_6244_0 = v_607_0 | v_26_0;
  assign v_6245_0 = v_6246_0 | v_8773_0;
  assign v_6246_0 = v_6247_0 | v_8772_0;
  assign v_6247_0 = v_589_0 ? v_6248_0 : 3'h0;
  assign v_6249_0 = v_6250_0 | v_6251_0;
  assign v_6250_0 = v_589_0 | v_601_0;
  assign v_6251_0 = v_607_0 | v_26_0;
  assign v_6252_0 = v_6253_0 | v_8769_0;
  assign v_6253_0 = v_6254_0 | v_8768_0;
  assign v_6254_0 = v_589_0 ? v_6255_0 : 3'h0;
  assign v_6256_0 = v_6257_0 | v_6258_0;
  assign v_6257_0 = v_589_0 | v_601_0;
  assign v_6258_0 = v_607_0 | v_26_0;
  assign v_6259_0 = v_6260_0 | v_8765_0;
  assign v_6260_0 = v_6261_0 | v_8764_0;
  assign v_6261_0 = v_589_0 ? v_6262_0 : 3'h0;
  assign v_6263_0 = v_6264_0 | v_6265_0;
  assign v_6264_0 = v_589_0 | v_601_0;
  assign v_6265_0 = v_607_0 | v_26_0;
  assign v_6266_0 = v_6267_0 | v_8761_0;
  assign v_6267_0 = v_6268_0 | v_8760_0;
  assign v_6268_0 = v_589_0 ? v_6269_0 : 3'h0;
  assign v_6270_0 = v_6271_0 | v_6272_0;
  assign v_6271_0 = v_589_0 | v_601_0;
  assign v_6272_0 = v_607_0 | v_26_0;
  assign v_6273_0 = v_6274_0 | v_8757_0;
  assign v_6274_0 = v_6275_0 | v_8756_0;
  assign v_6275_0 = v_589_0 ? v_6276_0 : 3'h0;
  assign v_6277_0 = v_6278_0 | v_6279_0;
  assign v_6278_0 = v_589_0 | v_601_0;
  assign v_6279_0 = v_607_0 | v_26_0;
  assign v_6280_0 = v_6281_0 | v_8753_0;
  assign v_6281_0 = v_6282_0 | v_8752_0;
  assign v_6282_0 = v_589_0 ? v_6283_0 : 3'h0;
  assign v_6284_0 = v_6285_0 | v_6286_0;
  assign v_6285_0 = v_589_0 | v_601_0;
  assign v_6286_0 = v_607_0 | v_26_0;
  assign v_6287_0 = v_6288_0 | v_8749_0;
  assign v_6288_0 = v_6289_0 | v_8748_0;
  assign v_6289_0 = v_589_0 ? v_6290_0 : 3'h0;
  assign v_6291_0 = v_6292_0 | v_6293_0;
  assign v_6292_0 = v_589_0 | v_601_0;
  assign v_6293_0 = v_607_0 | v_26_0;
  assign v_6294_0 = v_6295_0 | v_8745_0;
  assign v_6295_0 = v_6296_0 | v_8744_0;
  assign v_6296_0 = v_589_0 ? v_6297_0 : 3'h0;
  assign v_6298_0 = v_6299_0 | v_6300_0;
  assign v_6299_0 = v_589_0 | v_601_0;
  assign v_6300_0 = v_607_0 | v_26_0;
  assign v_6301_0 = v_6302_0 | v_8741_0;
  assign v_6302_0 = v_6303_0 | v_8740_0;
  assign v_6303_0 = v_589_0 ? v_6304_0 : 3'h0;
  assign v_6305_0 = v_6306_0 | v_6307_0;
  assign v_6306_0 = v_589_0 | v_601_0;
  assign v_6307_0 = v_607_0 | v_26_0;
  assign v_6308_0 = v_6309_0 | v_8737_0;
  assign v_6309_0 = v_6310_0 | v_8736_0;
  assign v_6310_0 = v_589_0 ? v_6311_0 : 3'h0;
  assign v_6312_0 = v_6313_0 | v_6314_0;
  assign v_6313_0 = v_589_0 | v_601_0;
  assign v_6314_0 = v_607_0 | v_26_0;
  assign v_6315_0 = v_6316_0 | v_8733_0;
  assign v_6316_0 = v_6317_0 | v_8732_0;
  assign v_6317_0 = v_589_0 ? v_6318_0 : 3'h0;
  assign v_6319_0 = v_6320_0 | v_6321_0;
  assign v_6320_0 = v_589_0 | v_601_0;
  assign v_6321_0 = v_607_0 | v_26_0;
  assign v_6322_0 = v_6323_0 | v_8729_0;
  assign v_6323_0 = v_6324_0 | v_8728_0;
  assign v_6324_0 = v_589_0 ? v_6325_0 : 3'h0;
  assign v_6326_0 = v_6327_0 | v_6328_0;
  assign v_6327_0 = v_589_0 | v_601_0;
  assign v_6328_0 = v_607_0 | v_26_0;
  assign v_6329_0 = v_6330_0 | v_8725_0;
  assign v_6330_0 = v_6331_0 | v_8724_0;
  assign v_6331_0 = v_589_0 ? v_6332_0 : 3'h0;
  assign v_6333_0 = v_6334_0 | v_6335_0;
  assign v_6334_0 = v_589_0 | v_601_0;
  assign v_6335_0 = v_607_0 | v_26_0;
  assign v_6336_0 = v_6337_0 | v_8721_0;
  assign v_6337_0 = v_6338_0 | v_8720_0;
  assign v_6338_0 = v_589_0 ? v_6339_0 : 3'h0;
  assign v_6340_0 = v_6341_0 | v_6342_0;
  assign v_6341_0 = v_589_0 | v_601_0;
  assign v_6342_0 = v_607_0 | v_26_0;
  assign v_6343_0 = v_6344_0 | v_8717_0;
  assign v_6344_0 = v_6345_0 | v_8716_0;
  assign v_6345_0 = v_589_0 ? v_6346_0 : 3'h0;
  assign v_6347_0 = v_6348_0 | v_6349_0;
  assign v_6348_0 = v_589_0 | v_601_0;
  assign v_6349_0 = v_607_0 | v_26_0;
  assign v_6350_0 = v_6351_0 | v_8713_0;
  assign v_6351_0 = v_6352_0 | v_8712_0;
  assign v_6352_0 = v_589_0 ? v_6353_0 : 3'h0;
  assign v_6354_0 = v_6355_0 | v_6356_0;
  assign v_6355_0 = v_589_0 | v_601_0;
  assign v_6356_0 = v_607_0 | v_26_0;
  assign v_6357_0 = v_6358_0 | v_8709_0;
  assign v_6358_0 = v_6359_0 | v_8708_0;
  assign v_6359_0 = v_589_0 ? v_6360_0 : 3'h0;
  assign v_6361_0 = v_6362_0 | v_6363_0;
  assign v_6362_0 = v_589_0 | v_601_0;
  assign v_6363_0 = v_607_0 | v_26_0;
  assign v_6364_0 = v_6365_0 | v_8705_0;
  assign v_6365_0 = v_6366_0 | v_8704_0;
  assign v_6366_0 = v_589_0 ? v_6367_0 : 3'h0;
  assign v_6368_0 = v_6369_0 | v_6370_0;
  assign v_6369_0 = v_589_0 | v_601_0;
  assign v_6370_0 = v_607_0 | v_26_0;
  assign v_6371_0 = v_6372_0 | v_8701_0;
  assign v_6372_0 = v_6373_0 | v_8700_0;
  assign v_6373_0 = v_589_0 ? v_6374_0 : 3'h0;
  assign v_6375_0 = v_6376_0 | v_6377_0;
  assign v_6376_0 = v_589_0 | v_601_0;
  assign v_6377_0 = v_607_0 | v_26_0;
  assign v_6378_0 = v_6379_0 | v_8697_0;
  assign v_6379_0 = v_6380_0 | v_8696_0;
  assign v_6380_0 = v_589_0 ? v_6381_0 : 3'h0;
  assign v_6382_0 = v_6383_0 | v_6384_0;
  assign v_6383_0 = v_589_0 | v_601_0;
  assign v_6384_0 = v_607_0 | v_26_0;
  assign v_6385_0 = v_6386_0 | v_8693_0;
  assign v_6386_0 = v_6387_0 | v_8692_0;
  assign v_6387_0 = v_589_0 ? v_6388_0 : 3'h0;
  assign v_6389_0 = v_6390_0 | v_6391_0;
  assign v_6390_0 = v_589_0 | v_601_0;
  assign v_6391_0 = v_607_0 | v_26_0;
  assign v_6392_0 = v_6393_0 | v_8689_0;
  assign v_6393_0 = v_6394_0 | v_8688_0;
  assign v_6394_0 = v_589_0 ? v_6395_0 : 3'h0;
  assign v_6396_0 = v_6397_0 | v_6398_0;
  assign v_6397_0 = v_589_0 | v_601_0;
  assign v_6398_0 = v_607_0 | v_26_0;
  assign v_6399_0 = v_6400_0 | v_8685_0;
  assign v_6400_0 = v_6401_0 | v_8684_0;
  assign v_6401_0 = v_589_0 ? v_6402_0 : 3'h0;
  assign v_6403_0 = v_6404_0 | v_6405_0;
  assign v_6404_0 = v_589_0 | v_601_0;
  assign v_6405_0 = v_607_0 | v_26_0;
  assign v_6406_0 = v_6407_0 | v_8681_0;
  assign v_6407_0 = v_6408_0 | v_8680_0;
  assign v_6408_0 = v_589_0 ? v_6409_0 : 3'h0;
  assign v_6410_0 = v_6411_0 | v_6412_0;
  assign v_6411_0 = v_589_0 | v_601_0;
  assign v_6412_0 = v_607_0 | v_26_0;
  assign v_6413_0 = v_6414_0 | v_8677_0;
  assign v_6414_0 = v_6415_0 | v_8676_0;
  assign v_6415_0 = v_589_0 ? v_6416_0 : 3'h0;
  assign v_6417_0 = v_6418_0 | v_6419_0;
  assign v_6418_0 = v_589_0 | v_601_0;
  assign v_6419_0 = v_607_0 | v_26_0;
  assign v_6420_0 = v_6421_0 | v_8673_0;
  assign v_6421_0 = v_6422_0 | v_8672_0;
  assign v_6422_0 = v_589_0 ? v_6423_0 : 3'h0;
  assign v_6424_0 = v_6425_0 | v_6426_0;
  assign v_6425_0 = v_589_0 | v_601_0;
  assign v_6426_0 = v_607_0 | v_26_0;
  assign v_6427_0 = v_6428_0 | v_8669_0;
  assign v_6428_0 = v_6429_0 | v_8668_0;
  assign v_6429_0 = v_589_0 ? v_6430_0 : 3'h0;
  assign v_6431_0 = v_6432_0 | v_6433_0;
  assign v_6432_0 = v_589_0 | v_601_0;
  assign v_6433_0 = v_607_0 | v_26_0;
  assign v_6434_0 = v_6435_0 | v_8665_0;
  assign v_6435_0 = v_6436_0 | v_8664_0;
  assign v_6436_0 = v_589_0 ? v_6437_0 : 3'h0;
  assign v_6438_0 = v_6439_0 | v_6440_0;
  assign v_6439_0 = v_589_0 | v_601_0;
  assign v_6440_0 = v_607_0 | v_26_0;
  assign v_6441_0 = v_6442_0 | v_8661_0;
  assign v_6442_0 = v_6443_0 | v_8660_0;
  assign v_6443_0 = v_589_0 ? v_6444_0 : 3'h0;
  assign v_6445_0 = v_6446_0 | v_6447_0;
  assign v_6446_0 = v_589_0 | v_601_0;
  assign v_6447_0 = v_607_0 | v_26_0;
  assign v_6448_0 = v_6449_0 | v_8657_0;
  assign v_6449_0 = v_6450_0 | v_8656_0;
  assign v_6450_0 = v_589_0 ? v_6451_0 : 3'h0;
  assign v_6452_0 = v_6453_0 | v_6454_0;
  assign v_6453_0 = v_589_0 | v_601_0;
  assign v_6454_0 = v_607_0 | v_26_0;
  assign v_6455_0 = v_6456_0 | v_8653_0;
  assign v_6456_0 = v_6457_0 | v_8652_0;
  assign v_6457_0 = v_589_0 ? v_6458_0 : 3'h0;
  assign v_6459_0 = v_6460_0 | v_6461_0;
  assign v_6460_0 = v_589_0 | v_601_0;
  assign v_6461_0 = v_607_0 | v_26_0;
  assign v_6462_0 = v_6463_0 | v_8649_0;
  assign v_6463_0 = v_6464_0 | v_8648_0;
  assign v_6464_0 = v_589_0 ? v_6465_0 : 3'h0;
  assign v_6466_0 = v_6467_0 | v_6468_0;
  assign v_6467_0 = v_589_0 | v_601_0;
  assign v_6468_0 = v_607_0 | v_26_0;
  assign v_6469_0 = v_6470_0 | v_8645_0;
  assign v_6470_0 = v_6471_0 | v_8644_0;
  assign v_6471_0 = v_589_0 ? v_6472_0 : 3'h0;
  assign v_6473_0 = v_6474_0 | v_6475_0;
  assign v_6474_0 = v_589_0 | v_601_0;
  assign v_6475_0 = v_607_0 | v_26_0;
  assign v_6476_0 = v_6477_0 | v_8641_0;
  assign v_6477_0 = v_6478_0 | v_8640_0;
  assign v_6478_0 = v_589_0 ? v_6479_0 : 3'h0;
  assign v_6480_0 = v_6481_0 | v_6482_0;
  assign v_6481_0 = v_589_0 | v_601_0;
  assign v_6482_0 = v_607_0 | v_26_0;
  assign v_6483_0 = v_6484_0 | v_8637_0;
  assign v_6484_0 = v_6485_0 | v_8636_0;
  assign v_6485_0 = v_589_0 ? v_6486_0 : 3'h0;
  assign v_6487_0 = v_6488_0 | v_6489_0;
  assign v_6488_0 = v_589_0 | v_601_0;
  assign v_6489_0 = v_607_0 | v_26_0;
  assign v_6490_0 = v_6491_0 | v_8633_0;
  assign v_6491_0 = v_6492_0 | v_8632_0;
  assign v_6492_0 = v_589_0 ? v_6493_0 : 3'h0;
  assign v_6494_0 = v_6495_0 | v_6496_0;
  assign v_6495_0 = v_589_0 | v_601_0;
  assign v_6496_0 = v_607_0 | v_26_0;
  assign v_6497_0 = v_6498_0 | v_8629_0;
  assign v_6498_0 = v_6499_0 | v_8628_0;
  assign v_6499_0 = v_589_0 ? v_6500_0 : 3'h0;
  assign v_6501_0 = v_6502_0 | v_6503_0;
  assign v_6502_0 = v_589_0 | v_601_0;
  assign v_6503_0 = v_607_0 | v_26_0;
  assign v_6504_0 = v_6505_0 | v_8625_0;
  assign v_6505_0 = v_6506_0 | v_8624_0;
  assign v_6506_0 = v_589_0 ? v_6507_0 : 3'h0;
  assign v_6508_0 = v_6509_0 | v_6510_0;
  assign v_6509_0 = v_589_0 | v_601_0;
  assign v_6510_0 = v_607_0 | v_26_0;
  assign v_6511_0 = v_6512_0 | v_8621_0;
  assign v_6512_0 = v_6513_0 | v_8620_0;
  assign v_6513_0 = v_589_0 ? v_6514_0 : 3'h0;
  assign v_6515_0 = v_6516_0 | v_6517_0;
  assign v_6516_0 = v_589_0 | v_601_0;
  assign v_6517_0 = v_607_0 | v_26_0;
  assign v_6518_0 = v_6519_0 | v_8617_0;
  assign v_6519_0 = v_6520_0 | v_8616_0;
  assign v_6520_0 = v_589_0 ? v_6521_0 : 3'h0;
  assign v_6522_0 = v_6523_0 | v_6524_0;
  assign v_6523_0 = v_589_0 | v_601_0;
  assign v_6524_0 = v_607_0 | v_26_0;
  assign v_6525_0 = v_6526_0 | v_8613_0;
  assign v_6526_0 = v_6527_0 | v_8612_0;
  assign v_6527_0 = v_589_0 ? v_6528_0 : 3'h0;
  assign v_6529_0 = v_6530_0 | v_6531_0;
  assign v_6530_0 = v_589_0 | v_601_0;
  assign v_6531_0 = v_607_0 | v_26_0;
  assign v_6532_0 = v_6533_0 | v_8609_0;
  assign v_6533_0 = v_6534_0 | v_8608_0;
  assign v_6534_0 = v_589_0 ? v_6535_0 : 3'h0;
  assign v_6536_0 = v_6537_0 | v_6538_0;
  assign v_6537_0 = v_589_0 | v_601_0;
  assign v_6538_0 = v_607_0 | v_26_0;
  assign v_6539_0 = v_6540_0 | v_8605_0;
  assign v_6540_0 = v_6541_0 | v_8604_0;
  assign v_6541_0 = v_589_0 ? v_6542_0 : 3'h0;
  assign v_6543_0 = v_6544_0 | v_6545_0;
  assign v_6544_0 = v_589_0 | v_601_0;
  assign v_6545_0 = v_607_0 | v_26_0;
  assign v_6546_0 = v_6547_0 | v_8601_0;
  assign v_6547_0 = v_6548_0 | v_8600_0;
  assign v_6548_0 = v_589_0 ? v_6549_0 : 3'h0;
  assign v_6550_0 = v_6551_0 | v_6552_0;
  assign v_6551_0 = v_589_0 | v_601_0;
  assign v_6552_0 = v_607_0 | v_26_0;
  assign v_6553_0 = v_6554_0 | v_8597_0;
  assign v_6554_0 = v_6555_0 | v_8596_0;
  assign v_6555_0 = v_589_0 ? v_6556_0 : 3'h0;
  assign v_6557_0 = v_6558_0 | v_6559_0;
  assign v_6558_0 = v_589_0 | v_601_0;
  assign v_6559_0 = v_607_0 | v_26_0;
  assign v_6560_0 = v_6561_0 | v_8593_0;
  assign v_6561_0 = v_6562_0 | v_8592_0;
  assign v_6562_0 = v_589_0 ? v_6563_0 : 3'h0;
  assign v_6564_0 = v_6565_0 | v_6566_0;
  assign v_6565_0 = v_589_0 | v_601_0;
  assign v_6566_0 = v_607_0 | v_26_0;
  assign v_6567_0 = v_6568_0 | v_8589_0;
  assign v_6568_0 = v_6569_0 | v_8588_0;
  assign v_6569_0 = v_589_0 ? v_6570_0 : 3'h0;
  assign v_6571_0 = v_6572_0 | v_6573_0;
  assign v_6572_0 = v_589_0 | v_601_0;
  assign v_6573_0 = v_607_0 | v_26_0;
  assign v_6574_0 = v_6575_0 | v_8585_0;
  assign v_6575_0 = v_6576_0 | v_8584_0;
  assign v_6576_0 = v_589_0 ? v_6577_0 : 3'h0;
  assign v_6578_0 = v_6579_0 | v_6580_0;
  assign v_6579_0 = v_589_0 | v_601_0;
  assign v_6580_0 = v_607_0 | v_26_0;
  assign v_6581_0 = v_6582_0 | v_8581_0;
  assign v_6582_0 = v_6583_0 | v_8580_0;
  assign v_6583_0 = v_589_0 ? v_6584_0 : 3'h0;
  assign v_6585_0 = v_6586_0 | v_6587_0;
  assign v_6586_0 = v_589_0 | v_601_0;
  assign v_6587_0 = v_607_0 | v_26_0;
  assign v_6588_0 = v_6589_0 | v_8577_0;
  assign v_6589_0 = v_6590_0 | v_8576_0;
  assign v_6590_0 = v_589_0 ? v_6591_0 : 3'h0;
  assign v_6592_0 = v_6593_0 | v_6594_0;
  assign v_6593_0 = v_589_0 | v_601_0;
  assign v_6594_0 = v_607_0 | v_26_0;
  assign v_6595_0 = v_6596_0 | v_8573_0;
  assign v_6596_0 = v_6597_0 | v_8572_0;
  assign v_6597_0 = v_589_0 ? v_6598_0 : 3'h0;
  assign v_6599_0 = v_6600_0 | v_6601_0;
  assign v_6600_0 = v_589_0 | v_601_0;
  assign v_6601_0 = v_607_0 | v_26_0;
  assign v_6602_0 = v_6603_0 | v_8569_0;
  assign v_6603_0 = v_6604_0 | v_8568_0;
  assign v_6604_0 = v_589_0 ? v_6605_0 : 3'h0;
  assign v_6606_0 = v_6607_0 | v_6608_0;
  assign v_6607_0 = v_589_0 | v_601_0;
  assign v_6608_0 = v_607_0 | v_26_0;
  assign v_6609_0 = v_6610_0 | v_8565_0;
  assign v_6610_0 = v_6611_0 | v_8564_0;
  assign v_6611_0 = v_589_0 ? v_6612_0 : 3'h0;
  assign v_6613_0 = v_6614_0 | v_6615_0;
  assign v_6614_0 = v_589_0 | v_601_0;
  assign v_6615_0 = v_607_0 | v_26_0;
  assign v_6616_0 = v_6617_0 | v_8561_0;
  assign v_6617_0 = v_6618_0 | v_8560_0;
  assign v_6618_0 = v_589_0 ? v_6619_0 : 3'h0;
  assign v_6620_0 = v_6621_0 | v_6622_0;
  assign v_6621_0 = v_589_0 | v_601_0;
  assign v_6622_0 = v_607_0 | v_26_0;
  assign v_6623_0 = v_6624_0 | v_8557_0;
  assign v_6624_0 = v_6625_0 | v_8556_0;
  assign v_6625_0 = v_589_0 ? v_6626_0 : 3'h0;
  assign v_6627_0 = v_6628_0 | v_6629_0;
  assign v_6628_0 = v_589_0 | v_601_0;
  assign v_6629_0 = v_607_0 | v_26_0;
  assign v_6630_0 = v_6631_0 | v_8553_0;
  assign v_6631_0 = v_6632_0 | v_8552_0;
  assign v_6632_0 = v_589_0 ? v_6633_0 : 3'h0;
  assign v_6634_0 = v_6635_0 | v_6636_0;
  assign v_6635_0 = v_589_0 | v_601_0;
  assign v_6636_0 = v_607_0 | v_26_0;
  assign v_6637_0 = v_6638_0 | v_8549_0;
  assign v_6638_0 = v_6639_0 | v_8548_0;
  assign v_6639_0 = v_589_0 ? v_6640_0 : 3'h0;
  assign v_6641_0 = v_6642_0 | v_6643_0;
  assign v_6642_0 = v_589_0 | v_601_0;
  assign v_6643_0 = v_607_0 | v_26_0;
  assign v_6644_0 = v_6645_0 | v_8545_0;
  assign v_6645_0 = v_6646_0 | v_8544_0;
  assign v_6646_0 = v_589_0 ? v_6647_0 : 3'h0;
  assign v_6648_0 = v_6649_0 | v_6650_0;
  assign v_6649_0 = v_589_0 | v_601_0;
  assign v_6650_0 = v_607_0 | v_26_0;
  assign v_6651_0 = v_6652_0 | v_8541_0;
  assign v_6652_0 = v_6653_0 | v_8540_0;
  assign v_6653_0 = v_589_0 ? v_6654_0 : 3'h0;
  assign v_6655_0 = v_6656_0 | v_6657_0;
  assign v_6656_0 = v_589_0 | v_601_0;
  assign v_6657_0 = v_607_0 | v_26_0;
  assign v_6658_0 = v_6659_0 | v_8537_0;
  assign v_6659_0 = v_6660_0 | v_8536_0;
  assign v_6660_0 = v_589_0 ? v_6661_0 : 3'h0;
  assign v_6662_0 = v_6663_0 | v_6664_0;
  assign v_6663_0 = v_589_0 | v_601_0;
  assign v_6664_0 = v_607_0 | v_26_0;
  assign v_6665_0 = v_6666_0 | v_8533_0;
  assign v_6666_0 = v_6667_0 | v_8532_0;
  assign v_6667_0 = v_589_0 ? v_6668_0 : 3'h0;
  assign v_6669_0 = v_6670_0 | v_6671_0;
  assign v_6670_0 = v_589_0 | v_601_0;
  assign v_6671_0 = v_607_0 | v_26_0;
  assign v_6672_0 = v_6673_0 | v_8529_0;
  assign v_6673_0 = v_6674_0 | v_8528_0;
  assign v_6674_0 = v_589_0 ? v_6675_0 : 3'h0;
  assign v_6676_0 = v_6677_0 | v_6678_0;
  assign v_6677_0 = v_589_0 | v_601_0;
  assign v_6678_0 = v_607_0 | v_26_0;
  assign v_6679_0 = v_6680_0 | v_8525_0;
  assign v_6680_0 = v_6681_0 | v_8524_0;
  assign v_6681_0 = v_589_0 ? v_6682_0 : 3'h0;
  assign v_6683_0 = v_6684_0 | v_6685_0;
  assign v_6684_0 = v_589_0 | v_601_0;
  assign v_6685_0 = v_607_0 | v_26_0;
  assign v_6686_0 = v_6687_0 | v_8521_0;
  assign v_6687_0 = v_6688_0 | v_8520_0;
  assign v_6688_0 = v_589_0 ? v_6689_0 : 3'h0;
  assign v_6690_0 = v_6691_0 | v_6692_0;
  assign v_6691_0 = v_589_0 | v_601_0;
  assign v_6692_0 = v_607_0 | v_26_0;
  assign v_6693_0 = v_6694_0 | v_8517_0;
  assign v_6694_0 = v_6695_0 | v_8516_0;
  assign v_6695_0 = v_589_0 ? v_6696_0 : 3'h0;
  assign v_6697_0 = v_6698_0 | v_6699_0;
  assign v_6698_0 = v_589_0 | v_601_0;
  assign v_6699_0 = v_607_0 | v_26_0;
  assign v_6700_0 = v_6701_0 | v_8513_0;
  assign v_6701_0 = v_6702_0 | v_8512_0;
  assign v_6702_0 = v_589_0 ? v_6703_0 : 3'h0;
  assign v_6704_0 = v_6705_0 | v_6706_0;
  assign v_6705_0 = v_589_0 | v_601_0;
  assign v_6706_0 = v_607_0 | v_26_0;
  assign v_6707_0 = v_6708_0 | v_8509_0;
  assign v_6708_0 = v_6709_0 | v_8508_0;
  assign v_6709_0 = v_589_0 ? v_6710_0 : 3'h0;
  assign v_6711_0 = v_6712_0 | v_6713_0;
  assign v_6712_0 = v_589_0 | v_601_0;
  assign v_6713_0 = v_607_0 | v_26_0;
  assign v_6714_0 = v_6715_0 | v_8505_0;
  assign v_6715_0 = v_6716_0 | v_8504_0;
  assign v_6716_0 = v_589_0 ? v_6717_0 : 3'h0;
  assign v_6718_0 = v_6719_0 | v_6720_0;
  assign v_6719_0 = v_589_0 | v_601_0;
  assign v_6720_0 = v_607_0 | v_26_0;
  assign v_6721_0 = v_6722_0 | v_8501_0;
  assign v_6722_0 = v_6723_0 | v_8500_0;
  assign v_6723_0 = v_589_0 ? v_6724_0 : 3'h0;
  assign v_6725_0 = v_6726_0 | v_6727_0;
  assign v_6726_0 = v_589_0 | v_601_0;
  assign v_6727_0 = v_607_0 | v_26_0;
  assign v_6728_0 = v_6729_0 | v_8497_0;
  assign v_6729_0 = v_6730_0 | v_8496_0;
  assign v_6730_0 = v_589_0 ? v_6731_0 : 3'h0;
  assign v_6732_0 = v_6733_0 | v_6734_0;
  assign v_6733_0 = v_589_0 | v_601_0;
  assign v_6734_0 = v_607_0 | v_26_0;
  assign v_6735_0 = v_6736_0 | v_8493_0;
  assign v_6736_0 = v_6737_0 | v_8492_0;
  assign v_6737_0 = v_589_0 ? v_6738_0 : 3'h0;
  assign v_6739_0 = v_6740_0 | v_6741_0;
  assign v_6740_0 = v_589_0 | v_601_0;
  assign v_6741_0 = v_607_0 | v_26_0;
  assign v_6742_0 = v_6743_0 | v_8489_0;
  assign v_6743_0 = v_6744_0 | v_8488_0;
  assign v_6744_0 = v_589_0 ? v_6745_0 : 3'h0;
  assign v_6746_0 = v_6747_0 | v_6748_0;
  assign v_6747_0 = v_589_0 | v_601_0;
  assign v_6748_0 = v_607_0 | v_26_0;
  assign v_6749_0 = v_6750_0 | v_8485_0;
  assign v_6750_0 = v_6751_0 | v_8484_0;
  assign v_6751_0 = v_589_0 ? v_6752_0 : 3'h0;
  assign v_6753_0 = v_6754_0 | v_6755_0;
  assign v_6754_0 = v_589_0 | v_601_0;
  assign v_6755_0 = v_607_0 | v_26_0;
  assign v_6756_0 = v_6757_0 | v_8481_0;
  assign v_6757_0 = v_6758_0 | v_8480_0;
  assign v_6758_0 = v_589_0 ? v_6759_0 : 3'h0;
  assign v_6760_0 = v_6761_0 | v_6762_0;
  assign v_6761_0 = v_589_0 | v_601_0;
  assign v_6762_0 = v_607_0 | v_26_0;
  assign v_6763_0 = v_6764_0 | v_8477_0;
  assign v_6764_0 = v_6765_0 | v_8476_0;
  assign v_6765_0 = v_589_0 ? v_6766_0 : 3'h0;
  assign v_6767_0 = v_6768_0 | v_6769_0;
  assign v_6768_0 = v_589_0 | v_601_0;
  assign v_6769_0 = v_607_0 | v_26_0;
  assign v_6770_0 = v_6771_0 | v_8473_0;
  assign v_6771_0 = v_6772_0 | v_8472_0;
  assign v_6772_0 = v_589_0 ? v_6773_0 : 3'h0;
  assign v_6774_0 = v_6775_0 | v_6776_0;
  assign v_6775_0 = v_589_0 | v_601_0;
  assign v_6776_0 = v_607_0 | v_26_0;
  assign v_6777_0 = v_6778_0 | v_8469_0;
  assign v_6778_0 = v_6779_0 | v_8468_0;
  assign v_6779_0 = v_589_0 ? v_6780_0 : 3'h0;
  assign v_6781_0 = v_6782_0 | v_6783_0;
  assign v_6782_0 = v_589_0 | v_601_0;
  assign v_6783_0 = v_607_0 | v_26_0;
  assign v_6784_0 = v_6785_0 | v_8465_0;
  assign v_6785_0 = v_6786_0 | v_8464_0;
  assign v_6786_0 = v_589_0 ? v_6787_0 : 3'h0;
  assign v_6788_0 = v_6789_0 | v_6790_0;
  assign v_6789_0 = v_589_0 | v_601_0;
  assign v_6790_0 = v_607_0 | v_26_0;
  assign v_6791_0 = v_6792_0 | v_8461_0;
  assign v_6792_0 = v_6793_0 | v_8460_0;
  assign v_6793_0 = v_589_0 ? v_6794_0 : 3'h0;
  assign v_6795_0 = v_6796_0 | v_6797_0;
  assign v_6796_0 = v_589_0 | v_601_0;
  assign v_6797_0 = v_607_0 | v_26_0;
  assign v_6798_0 = v_6799_0 | v_8457_0;
  assign v_6799_0 = v_6800_0 | v_8456_0;
  assign v_6800_0 = v_589_0 ? v_6801_0 : 3'h0;
  assign v_6802_0 = v_6803_0 | v_6804_0;
  assign v_6803_0 = v_589_0 | v_601_0;
  assign v_6804_0 = v_607_0 | v_26_0;
  assign v_6805_0 = v_6806_0 | v_8453_0;
  assign v_6806_0 = v_6807_0 | v_8452_0;
  assign v_6807_0 = v_589_0 ? v_6808_0 : 3'h0;
  assign v_6809_0 = v_6810_0 | v_6811_0;
  assign v_6810_0 = v_589_0 | v_601_0;
  assign v_6811_0 = v_607_0 | v_26_0;
  assign v_6812_0 = v_6813_0 | v_8449_0;
  assign v_6813_0 = v_6814_0 | v_8448_0;
  assign v_6814_0 = v_589_0 ? v_6815_0 : 3'h0;
  assign v_6816_0 = v_6817_0 | v_6818_0;
  assign v_6817_0 = v_589_0 | v_601_0;
  assign v_6818_0 = v_607_0 | v_26_0;
  assign v_6819_0 = v_6820_0 | v_8445_0;
  assign v_6820_0 = v_6821_0 | v_8444_0;
  assign v_6821_0 = v_589_0 ? v_6822_0 : 3'h0;
  assign v_6823_0 = v_6824_0 | v_6825_0;
  assign v_6824_0 = v_589_0 | v_601_0;
  assign v_6825_0 = v_607_0 | v_26_0;
  assign v_6826_0 = v_6827_0 | v_8441_0;
  assign v_6827_0 = v_6828_0 | v_8440_0;
  assign v_6828_0 = v_589_0 ? v_6829_0 : 3'h0;
  assign v_6830_0 = v_6831_0 | v_6832_0;
  assign v_6831_0 = v_589_0 | v_601_0;
  assign v_6832_0 = v_607_0 | v_26_0;
  assign v_6833_0 = v_6834_0 | v_8437_0;
  assign v_6834_0 = v_6835_0 | v_8436_0;
  assign v_6835_0 = v_589_0 ? v_6836_0 : 3'h0;
  assign v_6837_0 = v_6838_0 | v_6839_0;
  assign v_6838_0 = v_589_0 | v_601_0;
  assign v_6839_0 = v_607_0 | v_26_0;
  assign v_6840_0 = v_6841_0 | v_8433_0;
  assign v_6841_0 = v_6842_0 | v_8432_0;
  assign v_6842_0 = v_589_0 ? v_6843_0 : 3'h0;
  assign v_6844_0 = v_6845_0 | v_6846_0;
  assign v_6845_0 = v_589_0 | v_601_0;
  assign v_6846_0 = v_607_0 | v_26_0;
  assign v_6847_0 = v_6848_0 | v_8429_0;
  assign v_6848_0 = v_6849_0 | v_8428_0;
  assign v_6849_0 = v_589_0 ? v_6850_0 : 3'h0;
  assign v_6851_0 = v_6852_0 | v_6853_0;
  assign v_6852_0 = v_589_0 | v_601_0;
  assign v_6853_0 = v_607_0 | v_26_0;
  assign v_6854_0 = v_6855_0 | v_8425_0;
  assign v_6855_0 = v_6856_0 | v_8424_0;
  assign v_6856_0 = v_589_0 ? v_6857_0 : 3'h0;
  assign v_6858_0 = v_6859_0 | v_6860_0;
  assign v_6859_0 = v_589_0 | v_601_0;
  assign v_6860_0 = v_607_0 | v_26_0;
  assign v_6861_0 = v_6862_0 | v_8421_0;
  assign v_6862_0 = v_6863_0 | v_8420_0;
  assign v_6863_0 = v_589_0 ? v_6864_0 : 3'h0;
  assign v_6865_0 = v_6866_0 | v_6867_0;
  assign v_6866_0 = v_589_0 | v_601_0;
  assign v_6867_0 = v_607_0 | v_26_0;
  assign v_6868_0 = v_6869_0 | v_8417_0;
  assign v_6869_0 = v_6870_0 | v_8416_0;
  assign v_6870_0 = v_589_0 ? v_6871_0 : 3'h0;
  assign v_6872_0 = v_6873_0 | v_6874_0;
  assign v_6873_0 = v_589_0 | v_601_0;
  assign v_6874_0 = v_607_0 | v_26_0;
  assign v_6875_0 = v_6876_0 | v_8413_0;
  assign v_6876_0 = v_6877_0 | v_8412_0;
  assign v_6877_0 = v_589_0 ? v_6878_0 : 3'h0;
  assign v_6879_0 = v_6880_0 | v_6881_0;
  assign v_6880_0 = v_589_0 | v_601_0;
  assign v_6881_0 = v_607_0 | v_26_0;
  assign v_6882_0 = v_6883_0 | v_8409_0;
  assign v_6883_0 = v_6884_0 | v_8408_0;
  assign v_6884_0 = v_589_0 ? v_6885_0 : 3'h0;
  assign v_6886_0 = v_6887_0 | v_6888_0;
  assign v_6887_0 = v_589_0 | v_601_0;
  assign v_6888_0 = v_607_0 | v_26_0;
  assign v_6889_0 = v_6890_0 | v_8405_0;
  assign v_6890_0 = v_6891_0 | v_8404_0;
  assign v_6891_0 = v_589_0 ? v_6892_0 : 3'h0;
  assign v_6893_0 = v_6894_0 | v_6895_0;
  assign v_6894_0 = v_589_0 | v_601_0;
  assign v_6895_0 = v_607_0 | v_26_0;
  assign v_6896_0 = v_6897_0 | v_8401_0;
  assign v_6897_0 = v_6898_0 | v_8400_0;
  assign v_6898_0 = v_589_0 ? v_6899_0 : 3'h0;
  assign v_6900_0 = v_6901_0 | v_6902_0;
  assign v_6901_0 = v_589_0 | v_601_0;
  assign v_6902_0 = v_607_0 | v_26_0;
  assign v_6903_0 = v_6904_0 | v_8397_0;
  assign v_6904_0 = v_6905_0 | v_8396_0;
  assign v_6905_0 = v_589_0 ? v_6906_0 : 3'h0;
  assign v_6907_0 = v_6908_0 | v_6909_0;
  assign v_6908_0 = v_589_0 | v_601_0;
  assign v_6909_0 = v_607_0 | v_26_0;
  assign v_6910_0 = v_6911_0 | v_8393_0;
  assign v_6911_0 = v_6912_0 | v_8392_0;
  assign v_6912_0 = v_589_0 ? v_6913_0 : 3'h0;
  assign v_6914_0 = v_6915_0 | v_6916_0;
  assign v_6915_0 = v_589_0 | v_601_0;
  assign v_6916_0 = v_607_0 | v_26_0;
  assign v_6917_0 = v_6918_0 | v_8389_0;
  assign v_6918_0 = v_6919_0 | v_8388_0;
  assign v_6919_0 = v_589_0 ? v_6920_0 : 3'h0;
  assign v_6921_0 = v_6922_0 | v_6923_0;
  assign v_6922_0 = v_589_0 | v_601_0;
  assign v_6923_0 = v_607_0 | v_26_0;
  assign v_6924_0 = v_6925_0 | v_8385_0;
  assign v_6925_0 = v_6926_0 | v_8384_0;
  assign v_6926_0 = v_589_0 ? v_6927_0 : 3'h0;
  assign v_6928_0 = v_6929_0 | v_6930_0;
  assign v_6929_0 = v_589_0 | v_601_0;
  assign v_6930_0 = v_607_0 | v_26_0;
  assign v_6931_0 = v_6932_0 | v_8381_0;
  assign v_6932_0 = v_6933_0 | v_8380_0;
  assign v_6933_0 = v_589_0 ? v_6934_0 : 3'h0;
  assign v_6935_0 = v_6936_0 | v_6937_0;
  assign v_6936_0 = v_589_0 | v_601_0;
  assign v_6937_0 = v_607_0 | v_26_0;
  assign v_6938_0 = v_6939_0 | v_8377_0;
  assign v_6939_0 = v_6940_0 | v_8376_0;
  assign v_6940_0 = v_589_0 ? v_6941_0 : 3'h0;
  assign v_6942_0 = v_6943_0 | v_6944_0;
  assign v_6943_0 = v_589_0 | v_601_0;
  assign v_6944_0 = v_607_0 | v_26_0;
  assign v_6945_0 = v_6946_0 | v_8373_0;
  assign v_6946_0 = v_6947_0 | v_8372_0;
  assign v_6947_0 = v_589_0 ? v_6948_0 : 3'h0;
  assign v_6949_0 = v_6950_0 | v_6951_0;
  assign v_6950_0 = v_589_0 | v_601_0;
  assign v_6951_0 = v_607_0 | v_26_0;
  assign v_6952_0 = v_6953_0 | v_8369_0;
  assign v_6953_0 = v_6954_0 | v_8368_0;
  assign v_6954_0 = v_589_0 ? v_6955_0 : 3'h0;
  assign v_6956_0 = v_6957_0 | v_6958_0;
  assign v_6957_0 = v_589_0 | v_601_0;
  assign v_6958_0 = v_607_0 | v_26_0;
  assign v_6959_0 = v_6960_0 | v_8365_0;
  assign v_6960_0 = v_6961_0 | v_8364_0;
  assign v_6961_0 = v_589_0 ? v_6962_0 : 3'h0;
  assign v_6963_0 = v_6964_0 | v_6965_0;
  assign v_6964_0 = v_589_0 | v_601_0;
  assign v_6965_0 = v_607_0 | v_26_0;
  assign v_6966_0 = v_6967_0 | v_8361_0;
  assign v_6967_0 = v_6968_0 | v_8360_0;
  assign v_6968_0 = v_589_0 ? v_6969_0 : 3'h0;
  assign v_6970_0 = v_6971_0 | v_6972_0;
  assign v_6971_0 = v_589_0 | v_601_0;
  assign v_6972_0 = v_607_0 | v_26_0;
  assign v_6973_0 = v_6974_0 | v_8357_0;
  assign v_6974_0 = v_6975_0 | v_8356_0;
  assign v_6975_0 = v_589_0 ? v_6976_0 : 3'h0;
  assign v_6977_0 = v_6978_0 | v_6979_0;
  assign v_6978_0 = v_589_0 | v_601_0;
  assign v_6979_0 = v_607_0 | v_26_0;
  assign v_6980_0 = v_6981_0 | v_8353_0;
  assign v_6981_0 = v_6982_0 | v_8352_0;
  assign v_6982_0 = v_589_0 ? v_6983_0 : 3'h0;
  assign v_6984_0 = v_6985_0 | v_6986_0;
  assign v_6985_0 = v_589_0 | v_601_0;
  assign v_6986_0 = v_607_0 | v_26_0;
  assign v_6987_0 = v_6988_0 | v_8349_0;
  assign v_6988_0 = v_6989_0 | v_8348_0;
  assign v_6989_0 = v_589_0 ? v_6990_0 : 3'h0;
  assign v_6991_0 = v_6992_0 | v_6993_0;
  assign v_6992_0 = v_589_0 | v_601_0;
  assign v_6993_0 = v_607_0 | v_26_0;
  assign v_6994_0 = v_6995_0 | v_8345_0;
  assign v_6995_0 = v_6996_0 | v_8344_0;
  assign v_6996_0 = v_589_0 ? v_6997_0 : 3'h0;
  assign v_6998_0 = v_6999_0 | v_7000_0;
  assign v_6999_0 = v_589_0 | v_601_0;
  assign v_7000_0 = v_607_0 | v_26_0;
  assign v_7001_0 = v_7002_0 | v_8341_0;
  assign v_7002_0 = v_7003_0 | v_8340_0;
  assign v_7003_0 = v_589_0 ? v_7004_0 : 3'h0;
  assign v_7005_0 = v_7006_0 | v_7007_0;
  assign v_7006_0 = v_589_0 | v_601_0;
  assign v_7007_0 = v_607_0 | v_26_0;
  assign v_7008_0 = v_7009_0 | v_8337_0;
  assign v_7009_0 = v_7010_0 | v_8336_0;
  assign v_7010_0 = v_589_0 ? v_7011_0 : 3'h0;
  assign v_7012_0 = v_7013_0 | v_7014_0;
  assign v_7013_0 = v_589_0 | v_601_0;
  assign v_7014_0 = v_607_0 | v_26_0;
  assign v_7015_0 = v_7016_0 | v_8333_0;
  assign v_7016_0 = v_7017_0 | v_8332_0;
  assign v_7017_0 = v_589_0 ? v_7018_0 : 3'h0;
  assign v_7019_0 = v_7020_0 | v_7021_0;
  assign v_7020_0 = v_589_0 | v_601_0;
  assign v_7021_0 = v_607_0 | v_26_0;
  assign v_7022_0 = v_7023_0 | v_8329_0;
  assign v_7023_0 = v_7024_0 | v_8328_0;
  assign v_7024_0 = v_589_0 ? v_7025_0 : 3'h0;
  assign v_7026_0 = v_7027_0 | v_7028_0;
  assign v_7027_0 = v_589_0 | v_601_0;
  assign v_7028_0 = v_607_0 | v_26_0;
  assign v_7029_0 = v_7030_0 | v_8325_0;
  assign v_7030_0 = v_7031_0 | v_8324_0;
  assign v_7031_0 = v_589_0 ? v_7032_0 : 3'h0;
  assign v_7033_0 = v_7034_0 | v_7035_0;
  assign v_7034_0 = v_589_0 | v_601_0;
  assign v_7035_0 = v_607_0 | v_26_0;
  assign v_7036_0 = v_7037_0 | v_8321_0;
  assign v_7037_0 = v_7038_0 | v_8320_0;
  assign v_7038_0 = v_589_0 ? v_7039_0 : 3'h0;
  assign v_7040_0 = v_7041_0 | v_7042_0;
  assign v_7041_0 = v_589_0 | v_601_0;
  assign v_7042_0 = v_607_0 | v_26_0;
  assign v_7043_0 = v_7044_0 | v_8317_0;
  assign v_7044_0 = v_7045_0 | v_8316_0;
  assign v_7045_0 = v_589_0 ? v_7046_0 : 3'h0;
  assign v_7047_0 = v_7048_0 | v_7049_0;
  assign v_7048_0 = v_589_0 | v_601_0;
  assign v_7049_0 = v_607_0 | v_26_0;
  assign v_7050_0 = v_7051_0 | v_8313_0;
  assign v_7051_0 = v_7052_0 | v_8312_0;
  assign v_7052_0 = v_589_0 ? v_7053_0 : 3'h0;
  assign v_7054_0 = v_7055_0 | v_7056_0;
  assign v_7055_0 = v_589_0 | v_601_0;
  assign v_7056_0 = v_607_0 | v_26_0;
  assign v_7057_0 = v_7058_0 | v_8309_0;
  assign v_7058_0 = v_7059_0 | v_8308_0;
  assign v_7059_0 = v_589_0 ? v_7060_0 : 3'h0;
  assign v_7061_0 = v_7062_0 | v_7063_0;
  assign v_7062_0 = v_589_0 | v_601_0;
  assign v_7063_0 = v_607_0 | v_26_0;
  assign v_7064_0 = v_7065_0 | v_8305_0;
  assign v_7065_0 = v_7066_0 | v_8304_0;
  assign v_7066_0 = v_589_0 ? v_7067_0 : 3'h0;
  assign v_7068_0 = v_7069_0 | v_7070_0;
  assign v_7069_0 = v_589_0 | v_601_0;
  assign v_7070_0 = v_607_0 | v_26_0;
  assign v_7071_0 = v_7072_0 | v_8301_0;
  assign v_7072_0 = v_7073_0 | v_8300_0;
  assign v_7073_0 = v_589_0 ? v_7074_0 : 3'h0;
  assign v_7075_0 = v_7076_0 | v_7077_0;
  assign v_7076_0 = v_589_0 | v_601_0;
  assign v_7077_0 = v_607_0 | v_26_0;
  assign v_7078_0 = v_7079_0 | v_8297_0;
  assign v_7079_0 = v_7080_0 | v_8296_0;
  assign v_7080_0 = v_589_0 ? v_7081_0 : 3'h0;
  assign v_7082_0 = v_7083_0 | v_7084_0;
  assign v_7083_0 = v_589_0 | v_601_0;
  assign v_7084_0 = v_607_0 | v_26_0;
  assign v_7085_0 = v_7086_0 | v_8293_0;
  assign v_7086_0 = v_7087_0 | v_8292_0;
  assign v_7087_0 = v_589_0 ? v_7088_0 : 3'h0;
  assign v_7089_0 = v_7090_0 | v_7091_0;
  assign v_7090_0 = v_589_0 | v_601_0;
  assign v_7091_0 = v_607_0 | v_26_0;
  assign v_7092_0 = v_7093_0 | v_8289_0;
  assign v_7093_0 = v_7094_0 | v_8288_0;
  assign v_7094_0 = v_589_0 ? v_7095_0 : 3'h0;
  assign v_7096_0 = v_7097_0 | v_7098_0;
  assign v_7097_0 = v_589_0 | v_601_0;
  assign v_7098_0 = v_607_0 | v_26_0;
  assign v_7099_0 = v_7100_0 | v_8285_0;
  assign v_7100_0 = v_7101_0 | v_8284_0;
  assign v_7101_0 = v_589_0 ? v_7102_0 : 3'h0;
  assign v_7103_0 = v_7104_0 | v_7105_0;
  assign v_7104_0 = v_589_0 | v_601_0;
  assign v_7105_0 = v_607_0 | v_26_0;
  assign v_7106_0 = v_7107_0 | v_8281_0;
  assign v_7107_0 = v_7108_0 | v_8280_0;
  assign v_7108_0 = v_589_0 ? v_7109_0 : 3'h0;
  assign v_7110_0 = v_7111_0 | v_7112_0;
  assign v_7111_0 = v_589_0 | v_601_0;
  assign v_7112_0 = v_607_0 | v_26_0;
  assign v_7113_0 = v_7114_0 | v_8277_0;
  assign v_7114_0 = v_7115_0 | v_8276_0;
  assign v_7115_0 = v_589_0 ? v_7116_0 : 3'h0;
  assign v_7117_0 = v_7118_0 | v_7119_0;
  assign v_7118_0 = v_589_0 | v_601_0;
  assign v_7119_0 = v_607_0 | v_26_0;
  assign v_7120_0 = v_7121_0 | v_8273_0;
  assign v_7121_0 = v_7122_0 | v_8272_0;
  assign v_7122_0 = v_589_0 ? v_7123_0 : 3'h0;
  assign v_7124_0 = v_7125_0 | v_7126_0;
  assign v_7125_0 = v_589_0 | v_601_0;
  assign v_7126_0 = v_607_0 | v_26_0;
  assign v_7127_0 = v_7128_0 | v_8269_0;
  assign v_7128_0 = v_7129_0 | v_8268_0;
  assign v_7129_0 = v_589_0 ? v_7130_0 : 3'h0;
  assign v_7131_0 = v_7132_0 | v_7133_0;
  assign v_7132_0 = v_589_0 | v_601_0;
  assign v_7133_0 = v_607_0 | v_26_0;
  assign v_7134_0 = v_7135_0 | v_8265_0;
  assign v_7135_0 = v_7136_0 | v_8264_0;
  assign v_7136_0 = v_589_0 ? v_7137_0 : 3'h0;
  assign v_7138_0 = v_7139_0 | v_7140_0;
  assign v_7139_0 = v_589_0 | v_601_0;
  assign v_7140_0 = v_607_0 | v_26_0;
  assign v_7141_0 = v_7142_0 | v_8261_0;
  assign v_7142_0 = v_7143_0 | v_8260_0;
  assign v_7143_0 = v_589_0 ? v_7144_0 : 3'h0;
  assign v_7145_0 = v_7146_0 | v_7147_0;
  assign v_7146_0 = v_589_0 | v_601_0;
  assign v_7147_0 = v_607_0 | v_26_0;
  assign v_7148_0 = v_7149_0 | v_8257_0;
  assign v_7149_0 = v_7150_0 | v_8256_0;
  assign v_7150_0 = v_589_0 ? v_7151_0 : 3'h0;
  assign v_7152_0 = v_7153_0 | v_7154_0;
  assign v_7153_0 = v_589_0 | v_601_0;
  assign v_7154_0 = v_607_0 | v_26_0;
  assign v_7155_0 = v_7156_0 | v_8253_0;
  assign v_7156_0 = v_7157_0 | v_8252_0;
  assign v_7157_0 = v_589_0 ? v_7158_0 : 3'h0;
  assign v_7159_0 = v_7160_0 | v_7161_0;
  assign v_7160_0 = v_589_0 | v_601_0;
  assign v_7161_0 = v_607_0 | v_26_0;
  assign v_7162_0 = v_7163_0 | v_8249_0;
  assign v_7163_0 = v_7164_0 | v_8248_0;
  assign v_7164_0 = v_589_0 ? v_7165_0 : 3'h0;
  assign v_7166_0 = v_7167_0 | v_7168_0;
  assign v_7167_0 = v_589_0 | v_601_0;
  assign v_7168_0 = v_607_0 | v_26_0;
  assign v_7169_0 = v_7170_0 | v_8245_0;
  assign v_7170_0 = v_7171_0 | v_8244_0;
  assign v_7171_0 = v_589_0 ? v_7172_0 : 3'h0;
  assign v_7173_0 = v_7174_0 | v_7175_0;
  assign v_7174_0 = v_589_0 | v_601_0;
  assign v_7175_0 = v_607_0 | v_26_0;
  assign v_7176_0 = v_7177_0 | v_8241_0;
  assign v_7177_0 = v_7178_0 | v_8240_0;
  assign v_7178_0 = v_589_0 ? v_7179_0 : 3'h0;
  assign v_7180_0 = v_7181_0 | v_7182_0;
  assign v_7181_0 = v_589_0 | v_601_0;
  assign v_7182_0 = v_607_0 | v_26_0;
  assign v_7183_0 = v_7184_0 | v_8237_0;
  assign v_7184_0 = v_7185_0 | v_8236_0;
  assign v_7185_0 = v_589_0 ? v_7186_0 : 3'h0;
  assign v_7187_0 = v_7188_0 | v_7189_0;
  assign v_7188_0 = v_589_0 | v_601_0;
  assign v_7189_0 = v_607_0 | v_26_0;
  assign v_7190_0 = v_7191_0 | v_8233_0;
  assign v_7191_0 = v_7192_0 | v_8232_0;
  assign v_7192_0 = v_589_0 ? v_7193_0 : 3'h0;
  assign v_7194_0 = v_7195_0 | v_7196_0;
  assign v_7195_0 = v_589_0 | v_601_0;
  assign v_7196_0 = v_607_0 | v_26_0;
  assign v_7197_0 = v_7198_0 | v_8229_0;
  assign v_7198_0 = v_7199_0 | v_8228_0;
  assign v_7199_0 = v_589_0 ? v_7200_0 : 3'h0;
  assign v_7201_0 = v_7202_0 | v_7203_0;
  assign v_7202_0 = v_589_0 | v_601_0;
  assign v_7203_0 = v_607_0 | v_26_0;
  assign v_7204_0 = v_7205_0 | v_8225_0;
  assign v_7205_0 = v_7206_0 | v_8224_0;
  assign v_7206_0 = v_589_0 ? v_7207_0 : 3'h0;
  assign v_7208_0 = v_7209_0 | v_7210_0;
  assign v_7209_0 = v_589_0 | v_601_0;
  assign v_7210_0 = v_607_0 | v_26_0;
  assign v_7211_0 = v_7212_0 | v_8221_0;
  assign v_7212_0 = v_7213_0 | v_8220_0;
  assign v_7213_0 = v_589_0 ? v_7214_0 : 3'h0;
  assign v_7215_0 = v_7216_0 | v_7217_0;
  assign v_7216_0 = v_589_0 | v_601_0;
  assign v_7217_0 = v_607_0 | v_26_0;
  assign v_7218_0 = v_7219_0 | v_8217_0;
  assign v_7219_0 = v_7220_0 | v_8216_0;
  assign v_7220_0 = v_589_0 ? v_7221_0 : 3'h0;
  assign v_7222_0 = v_7223_0 | v_7224_0;
  assign v_7223_0 = v_589_0 | v_601_0;
  assign v_7224_0 = v_607_0 | v_26_0;
  assign v_7225_0 = v_7226_0 | v_8213_0;
  assign v_7226_0 = v_7227_0 | v_8212_0;
  assign v_7227_0 = v_589_0 ? v_7228_0 : 3'h0;
  assign v_7229_0 = v_7230_0 | v_7231_0;
  assign v_7230_0 = v_589_0 | v_601_0;
  assign v_7231_0 = v_607_0 | v_26_0;
  assign v_7232_0 = v_7233_0 | v_8209_0;
  assign v_7233_0 = v_7234_0 | v_8208_0;
  assign v_7234_0 = v_589_0 ? v_7235_0 : 3'h0;
  assign v_7236_0 = v_7237_0 | v_7238_0;
  assign v_7237_0 = v_589_0 | v_601_0;
  assign v_7238_0 = v_607_0 | v_26_0;
  assign v_7239_0 = v_7240_0 | v_8205_0;
  assign v_7240_0 = v_7241_0 | v_8204_0;
  assign v_7241_0 = v_589_0 ? v_7242_0 : 3'h0;
  assign v_7243_0 = v_7244_0 | v_7245_0;
  assign v_7244_0 = v_589_0 | v_601_0;
  assign v_7245_0 = v_607_0 | v_26_0;
  assign v_7246_0 = v_7247_0 | v_8201_0;
  assign v_7247_0 = v_7248_0 | v_8200_0;
  assign v_7248_0 = v_589_0 ? v_7249_0 : 3'h0;
  assign v_7250_0 = v_7251_0 | v_7252_0;
  assign v_7251_0 = v_589_0 | v_601_0;
  assign v_7252_0 = v_607_0 | v_26_0;
  assign v_7253_0 = v_7254_0 | v_8197_0;
  assign v_7254_0 = v_7255_0 | v_8196_0;
  assign v_7255_0 = v_589_0 ? v_7256_0 : 3'h0;
  assign v_7257_0 = v_7258_0 | v_7259_0;
  assign v_7258_0 = v_589_0 | v_601_0;
  assign v_7259_0 = v_607_0 | v_26_0;
  assign v_7260_0 = v_7261_0 | v_8193_0;
  assign v_7261_0 = v_7262_0 | v_8192_0;
  assign v_7262_0 = v_589_0 ? v_7263_0 : 3'h0;
  assign v_7264_0 = v_7265_0 | v_7266_0;
  assign v_7265_0 = v_589_0 | v_601_0;
  assign v_7266_0 = v_607_0 | v_26_0;
  assign v_7267_0 = v_7268_0 | v_8189_0;
  assign v_7268_0 = v_7269_0 | v_8188_0;
  assign v_7269_0 = v_589_0 ? v_7270_0 : 3'h0;
  assign v_7271_0 = v_7272_0 | v_7273_0;
  assign v_7272_0 = v_589_0 | v_601_0;
  assign v_7273_0 = v_607_0 | v_26_0;
  assign v_7274_0 = v_7275_0 | v_8185_0;
  assign v_7275_0 = v_7276_0 | v_8184_0;
  assign v_7276_0 = v_589_0 ? v_7277_0 : 3'h0;
  assign v_7278_0 = v_7279_0 | v_7280_0;
  assign v_7279_0 = v_589_0 | v_601_0;
  assign v_7280_0 = v_607_0 | v_26_0;
  assign v_7281_0 = v_7282_0 | v_8181_0;
  assign v_7282_0 = v_7283_0 | v_8180_0;
  assign v_7283_0 = v_589_0 ? v_7284_0 : 3'h0;
  assign v_7285_0 = v_7286_0 | v_7287_0;
  assign v_7286_0 = v_589_0 | v_601_0;
  assign v_7287_0 = v_607_0 | v_26_0;
  assign v_7288_0 = v_7289_0 | v_8177_0;
  assign v_7289_0 = v_7290_0 | v_8176_0;
  assign v_7290_0 = v_589_0 ? v_7291_0 : 3'h0;
  assign v_7292_0 = v_7293_0 | v_7294_0;
  assign v_7293_0 = v_589_0 | v_601_0;
  assign v_7294_0 = v_607_0 | v_26_0;
  assign v_7295_0 = v_7296_0 | v_8173_0;
  assign v_7296_0 = v_7297_0 | v_8172_0;
  assign v_7297_0 = v_589_0 ? v_7298_0 : 3'h0;
  assign v_7299_0 = v_7300_0 | v_7301_0;
  assign v_7300_0 = v_589_0 | v_601_0;
  assign v_7301_0 = v_607_0 | v_26_0;
  assign v_7302_0 = v_7303_0 | v_8169_0;
  assign v_7303_0 = v_7304_0 | v_8168_0;
  assign v_7304_0 = v_589_0 ? v_7305_0 : 3'h0;
  assign v_7306_0 = v_7307_0 | v_7308_0;
  assign v_7307_0 = v_589_0 | v_601_0;
  assign v_7308_0 = v_607_0 | v_26_0;
  assign v_7309_0 = v_7310_0 | v_8165_0;
  assign v_7310_0 = v_7311_0 | v_8164_0;
  assign v_7311_0 = v_589_0 ? v_7312_0 : 3'h0;
  assign v_7313_0 = v_7314_0 | v_7315_0;
  assign v_7314_0 = v_589_0 | v_601_0;
  assign v_7315_0 = v_607_0 | v_26_0;
  assign v_7316_0 = v_7317_0 | v_8161_0;
  assign v_7317_0 = v_7318_0 | v_8160_0;
  assign v_7318_0 = v_589_0 ? v_7319_0 : 3'h0;
  assign v_7320_0 = v_7321_0 | v_7322_0;
  assign v_7321_0 = v_589_0 | v_601_0;
  assign v_7322_0 = v_607_0 | v_26_0;
  assign v_7323_0 = v_7324_0 | v_8157_0;
  assign v_7324_0 = v_7325_0 | v_8156_0;
  assign v_7325_0 = v_589_0 ? v_7326_0 : 3'h0;
  assign v_7327_0 = v_7328_0 | v_7329_0;
  assign v_7328_0 = v_589_0 | v_601_0;
  assign v_7329_0 = v_607_0 | v_26_0;
  assign v_7330_0 = v_7331_0 | v_8153_0;
  assign v_7331_0 = v_7332_0 | v_8152_0;
  assign v_7332_0 = v_589_0 ? v_7333_0 : 3'h0;
  assign v_7334_0 = v_7335_0 | v_7336_0;
  assign v_7335_0 = v_589_0 | v_601_0;
  assign v_7336_0 = v_607_0 | v_26_0;
  assign v_7337_0 = v_7338_0 | v_8149_0;
  assign v_7338_0 = v_7339_0 | v_8148_0;
  assign v_7339_0 = v_589_0 ? v_7340_0 : 3'h0;
  assign v_7341_0 = v_7342_0 | v_7343_0;
  assign v_7342_0 = v_589_0 | v_601_0;
  assign v_7343_0 = v_607_0 | v_26_0;
  assign v_7344_0 = v_7345_0 | v_8145_0;
  assign v_7345_0 = v_7346_0 | v_8144_0;
  assign v_7346_0 = v_589_0 ? v_7347_0 : 3'h0;
  assign v_7348_0 = v_7349_0 | v_7350_0;
  assign v_7349_0 = v_589_0 | v_601_0;
  assign v_7350_0 = v_607_0 | v_26_0;
  assign v_7351_0 = v_7352_0 | v_8141_0;
  assign v_7352_0 = v_7353_0 | v_8140_0;
  assign v_7353_0 = v_589_0 ? v_7354_0 : 3'h0;
  assign v_7355_0 = v_7356_0 | v_7357_0;
  assign v_7356_0 = v_589_0 | v_601_0;
  assign v_7357_0 = v_607_0 | v_26_0;
  assign v_7358_0 = v_7359_0 | v_8137_0;
  assign v_7359_0 = v_7360_0 | v_8136_0;
  assign v_7360_0 = v_589_0 ? v_7361_0 : 3'h0;
  assign v_7362_0 = v_7363_0 | v_7364_0;
  assign v_7363_0 = v_589_0 | v_601_0;
  assign v_7364_0 = v_607_0 | v_26_0;
  assign v_7365_0 = v_7366_0 | v_8133_0;
  assign v_7366_0 = v_7367_0 | v_8132_0;
  assign v_7367_0 = v_589_0 ? v_7368_0 : 3'h0;
  assign v_7369_0 = v_7370_0 | v_7371_0;
  assign v_7370_0 = v_589_0 | v_601_0;
  assign v_7371_0 = v_607_0 | v_26_0;
  assign v_7372_0 = v_7373_0 | v_8129_0;
  assign v_7373_0 = v_7374_0 | v_8128_0;
  assign v_7374_0 = v_589_0 ? v_7375_0 : 3'h0;
  assign v_7376_0 = v_7377_0 | v_7378_0;
  assign v_7377_0 = v_589_0 | v_601_0;
  assign v_7378_0 = v_607_0 | v_26_0;
  assign v_7379_0 = v_7380_0 | v_8125_0;
  assign v_7380_0 = v_7381_0 | v_8124_0;
  assign v_7381_0 = v_589_0 ? v_7382_0 : 3'h0;
  assign v_7383_0 = v_7384_0 | v_7385_0;
  assign v_7384_0 = v_589_0 | v_601_0;
  assign v_7385_0 = v_607_0 | v_26_0;
  assign v_7386_0 = v_7387_0 | v_8121_0;
  assign v_7387_0 = v_7388_0 | v_8120_0;
  assign v_7388_0 = v_589_0 ? v_7389_0 : 3'h0;
  assign v_7390_0 = v_7391_0 | v_7392_0;
  assign v_7391_0 = v_589_0 | v_601_0;
  assign v_7392_0 = v_607_0 | v_26_0;
  assign v_7393_0 = v_7394_0 | v_8117_0;
  assign v_7394_0 = v_7395_0 | v_8116_0;
  assign v_7395_0 = v_589_0 ? v_7396_0 : 3'h0;
  assign v_7397_0 = v_7398_0 | v_7399_0;
  assign v_7398_0 = v_589_0 | v_601_0;
  assign v_7399_0 = v_607_0 | v_26_0;
  assign v_7400_0 = v_7401_0 | v_8113_0;
  assign v_7401_0 = v_7402_0 | v_8112_0;
  assign v_7402_0 = v_589_0 ? v_7403_0 : 3'h0;
  assign v_7404_0 = v_7405_0 | v_7406_0;
  assign v_7405_0 = v_589_0 | v_601_0;
  assign v_7406_0 = v_607_0 | v_26_0;
  assign v_7407_0 = v_7408_0 | v_8109_0;
  assign v_7408_0 = v_7409_0 | v_8108_0;
  assign v_7409_0 = v_589_0 ? v_7410_0 : 3'h0;
  assign v_7411_0 = v_7412_0 | v_7413_0;
  assign v_7412_0 = v_589_0 | v_601_0;
  assign v_7413_0 = v_607_0 | v_26_0;
  assign v_7414_0 = v_7415_0 | v_8105_0;
  assign v_7415_0 = v_7416_0 | v_8104_0;
  assign v_7416_0 = v_589_0 ? v_7417_0 : 3'h0;
  assign v_7418_0 = v_7419_0 | v_7420_0;
  assign v_7419_0 = v_589_0 | v_601_0;
  assign v_7420_0 = v_607_0 | v_26_0;
  assign v_7421_0 = v_7422_0 | v_8101_0;
  assign v_7422_0 = v_7423_0 | v_8100_0;
  assign v_7423_0 = v_589_0 ? v_7424_0 : 3'h0;
  assign v_7425_0 = v_7426_0 | v_7427_0;
  assign v_7426_0 = v_589_0 | v_601_0;
  assign v_7427_0 = v_607_0 | v_26_0;
  assign v_7428_0 = v_7429_0 | v_8097_0;
  assign v_7429_0 = v_7430_0 | v_8096_0;
  assign v_7430_0 = v_589_0 ? v_7431_0 : 3'h0;
  assign v_7432_0 = v_7433_0 | v_7434_0;
  assign v_7433_0 = v_589_0 | v_601_0;
  assign v_7434_0 = v_607_0 | v_26_0;
  assign v_7435_0 = v_7436_0 | v_8093_0;
  assign v_7436_0 = v_7437_0 | v_8092_0;
  assign v_7437_0 = v_589_0 ? v_7438_0 : 3'h0;
  assign v_7439_0 = v_7440_0 | v_7441_0;
  assign v_7440_0 = v_589_0 | v_601_0;
  assign v_7441_0 = v_607_0 | v_26_0;
  assign v_7442_0 = v_7443_0 | v_8089_0;
  assign v_7443_0 = v_7444_0 | v_8088_0;
  assign v_7444_0 = v_589_0 ? v_7445_0 : 3'h0;
  assign v_7446_0 = v_7447_0 | v_7448_0;
  assign v_7447_0 = v_589_0 | v_601_0;
  assign v_7448_0 = v_607_0 | v_26_0;
  assign v_7449_0 = v_7450_0 | v_8085_0;
  assign v_7450_0 = v_7451_0 | v_8084_0;
  assign v_7451_0 = v_589_0 ? v_7452_0 : 3'h0;
  assign v_7453_0 = v_7454_0 | v_7455_0;
  assign v_7454_0 = v_589_0 | v_601_0;
  assign v_7455_0 = v_607_0 | v_26_0;
  assign v_7456_0 = v_7457_0 | v_8081_0;
  assign v_7457_0 = v_7458_0 | v_8080_0;
  assign v_7458_0 = v_589_0 ? v_7459_0 : 3'h0;
  assign v_7460_0 = v_7461_0 | v_7462_0;
  assign v_7461_0 = v_589_0 | v_601_0;
  assign v_7462_0 = v_607_0 | v_26_0;
  assign v_7463_0 = v_7464_0 | v_8077_0;
  assign v_7464_0 = v_7465_0 | v_8076_0;
  assign v_7465_0 = v_589_0 ? v_7466_0 : 3'h0;
  assign v_7467_0 = v_7468_0 | v_7469_0;
  assign v_7468_0 = v_589_0 | v_601_0;
  assign v_7469_0 = v_607_0 | v_26_0;
  assign v_7470_0 = v_7471_0 | v_8073_0;
  assign v_7471_0 = v_7472_0 | v_8072_0;
  assign v_7472_0 = v_589_0 ? v_7473_0 : 3'h0;
  assign v_7474_0 = v_7475_0 | v_7476_0;
  assign v_7475_0 = v_589_0 | v_601_0;
  assign v_7476_0 = v_607_0 | v_26_0;
  assign v_7477_0 = v_7478_0 | v_8069_0;
  assign v_7478_0 = v_7479_0 | v_8068_0;
  assign v_7479_0 = v_589_0 ? v_7480_0 : 3'h0;
  assign v_7481_0 = v_7482_0 | v_7483_0;
  assign v_7482_0 = v_589_0 | v_601_0;
  assign v_7483_0 = v_607_0 | v_26_0;
  assign v_7484_0 = v_7485_0 | v_8065_0;
  assign v_7485_0 = v_7486_0 | v_8064_0;
  assign v_7486_0 = v_589_0 ? v_7487_0 : 3'h0;
  assign v_7488_0 = v_7489_0 | v_7490_0;
  assign v_7489_0 = v_589_0 | v_601_0;
  assign v_7490_0 = v_607_0 | v_26_0;
  assign v_7491_0 = v_7492_0 | v_8061_0;
  assign v_7492_0 = v_7493_0 | v_8060_0;
  assign v_7493_0 = v_589_0 ? v_7494_0 : 3'h0;
  assign v_7495_0 = v_7496_0 | v_7497_0;
  assign v_7496_0 = v_589_0 | v_601_0;
  assign v_7497_0 = v_607_0 | v_26_0;
  assign v_7498_0 = v_7499_0 | v_8057_0;
  assign v_7499_0 = v_7500_0 | v_8056_0;
  assign v_7500_0 = v_589_0 ? v_7501_0 : 3'h0;
  assign v_7502_0 = v_7503_0 | v_7504_0;
  assign v_7503_0 = v_589_0 | v_601_0;
  assign v_7504_0 = v_607_0 | v_26_0;
  assign v_7505_0 = v_7506_0 | v_8053_0;
  assign v_7506_0 = v_7507_0 | v_8052_0;
  assign v_7507_0 = v_589_0 ? v_7508_0 : 3'h0;
  assign v_7509_0 = v_7510_0 | v_7511_0;
  assign v_7510_0 = v_589_0 | v_601_0;
  assign v_7511_0 = v_607_0 | v_26_0;
  assign v_7512_0 = v_7513_0 | v_8049_0;
  assign v_7513_0 = v_7514_0 | v_8048_0;
  assign v_7514_0 = v_589_0 ? v_7515_0 : 3'h0;
  assign v_7516_0 = v_7517_0 | v_7518_0;
  assign v_7517_0 = v_589_0 | v_601_0;
  assign v_7518_0 = v_607_0 | v_26_0;
  assign v_7519_0 = v_7520_0 | v_8045_0;
  assign v_7520_0 = v_7521_0 | v_8044_0;
  assign v_7521_0 = v_589_0 ? v_7522_0 : 3'h0;
  assign v_7523_0 = v_7524_0 | v_7525_0;
  assign v_7524_0 = v_589_0 | v_601_0;
  assign v_7525_0 = v_607_0 | v_26_0;
  assign v_7526_0 = v_7527_0 | v_8041_0;
  assign v_7527_0 = v_7528_0 | v_8040_0;
  assign v_7528_0 = v_589_0 ? v_7529_0 : 3'h0;
  assign v_7530_0 = v_7531_0 | v_7532_0;
  assign v_7531_0 = v_589_0 | v_601_0;
  assign v_7532_0 = v_607_0 | v_26_0;
  assign v_7533_0 = v_7534_0 | v_8037_0;
  assign v_7534_0 = v_7535_0 | v_8036_0;
  assign v_7535_0 = v_589_0 ? v_7536_0 : 3'h0;
  assign v_7537_0 = v_7538_0 | v_7539_0;
  assign v_7538_0 = v_589_0 | v_601_0;
  assign v_7539_0 = v_607_0 | v_26_0;
  assign v_7540_0 = v_7541_0 | v_8033_0;
  assign v_7541_0 = v_7542_0 | v_8032_0;
  assign v_7542_0 = v_589_0 ? v_7543_0 : 3'h0;
  assign v_7544_0 = v_7545_0 | v_7546_0;
  assign v_7545_0 = v_589_0 | v_601_0;
  assign v_7546_0 = v_607_0 | v_26_0;
  assign v_7547_0 = v_7548_0 | v_8029_0;
  assign v_7548_0 = v_7549_0 | v_8028_0;
  assign v_7549_0 = v_589_0 ? v_7550_0 : 3'h0;
  assign v_7551_0 = v_7552_0 | v_7553_0;
  assign v_7552_0 = v_589_0 | v_601_0;
  assign v_7553_0 = v_607_0 | v_26_0;
  assign v_7554_0 = v_7555_0 | v_8025_0;
  assign v_7555_0 = v_7556_0 | v_8024_0;
  assign v_7556_0 = v_589_0 ? v_7557_0 : 3'h0;
  assign v_7558_0 = v_7559_0 | v_7560_0;
  assign v_7559_0 = v_589_0 | v_601_0;
  assign v_7560_0 = v_607_0 | v_26_0;
  assign v_7561_0 = v_7562_0 | v_8021_0;
  assign v_7562_0 = v_7563_0 | v_8020_0;
  assign v_7563_0 = v_589_0 ? v_7564_0 : 3'h0;
  assign v_7565_0 = v_7566_0 | v_7567_0;
  assign v_7566_0 = v_589_0 | v_601_0;
  assign v_7567_0 = v_607_0 | v_26_0;
  assign v_7568_0 = v_7569_0 | v_8017_0;
  assign v_7569_0 = v_7570_0 | v_8016_0;
  assign v_7570_0 = v_589_0 ? v_7571_0 : 3'h0;
  assign v_7572_0 = v_7573_0 | v_7574_0;
  assign v_7573_0 = v_589_0 | v_601_0;
  assign v_7574_0 = v_607_0 | v_26_0;
  assign v_7575_0 = v_7576_0 | v_8013_0;
  assign v_7576_0 = v_7577_0 | v_8012_0;
  assign v_7577_0 = v_589_0 ? v_7578_0 : 3'h0;
  assign v_7579_0 = v_7580_0 | v_7581_0;
  assign v_7580_0 = v_589_0 | v_601_0;
  assign v_7581_0 = v_607_0 | v_26_0;
  assign v_7582_0 = v_7583_0 | v_8009_0;
  assign v_7583_0 = v_7584_0 | v_8008_0;
  assign v_7584_0 = v_589_0 ? v_7585_0 : 3'h0;
  assign v_7586_0 = v_7587_0 | v_7588_0;
  assign v_7587_0 = v_589_0 | v_601_0;
  assign v_7588_0 = v_607_0 | v_26_0;
  assign v_7589_0 = v_7590_0 | v_8005_0;
  assign v_7590_0 = v_7591_0 | v_8004_0;
  assign v_7591_0 = v_589_0 ? v_7592_0 : 3'h0;
  assign v_7593_0 = v_7594_0 | v_7595_0;
  assign v_7594_0 = v_589_0 | v_601_0;
  assign v_7595_0 = v_607_0 | v_26_0;
  assign v_7596_0 = v_7597_0 | v_8001_0;
  assign v_7597_0 = v_7598_0 | v_8000_0;
  assign v_7598_0 = v_589_0 ? v_7599_0 : 3'h0;
  assign v_7600_0 = v_7601_0 | v_7602_0;
  assign v_7601_0 = v_589_0 | v_601_0;
  assign v_7602_0 = v_607_0 | v_26_0;
  assign v_7603_0 = v_7604_0 | v_7997_0;
  assign v_7604_0 = v_7605_0 | v_7996_0;
  assign v_7605_0 = v_589_0 ? v_7606_0 : 3'h0;
  assign v_7607_0 = v_7608_0 | v_7609_0;
  assign v_7608_0 = v_589_0 | v_601_0;
  assign v_7609_0 = v_607_0 | v_26_0;
  assign v_7610_0 = v_7611_0 | v_7993_0;
  assign v_7611_0 = v_7612_0 | v_7992_0;
  assign v_7612_0 = v_589_0 ? v_7613_0 : 3'h0;
  assign v_7614_0 = v_7615_0 | v_7616_0;
  assign v_7615_0 = v_589_0 | v_601_0;
  assign v_7616_0 = v_607_0 | v_26_0;
  assign v_7617_0 = v_7618_0 | v_7989_0;
  assign v_7618_0 = v_7619_0 | v_7988_0;
  assign v_7619_0 = v_589_0 ? v_7620_0 : 3'h0;
  assign v_7621_0 = v_7622_0 | v_7623_0;
  assign v_7622_0 = v_589_0 | v_601_0;
  assign v_7623_0 = v_607_0 | v_26_0;
  assign v_7624_0 = v_7625_0 | v_7985_0;
  assign v_7625_0 = v_7626_0 | v_7984_0;
  assign v_7626_0 = v_589_0 ? v_7627_0 : 3'h0;
  assign v_7628_0 = v_7629_0 | v_7630_0;
  assign v_7629_0 = v_589_0 | v_601_0;
  assign v_7630_0 = v_607_0 | v_26_0;
  assign v_7631_0 = v_7632_0 | v_7981_0;
  assign v_7632_0 = v_7633_0 | v_7980_0;
  assign v_7633_0 = v_589_0 ? v_7634_0 : 3'h0;
  assign v_7635_0 = v_7636_0 | v_7637_0;
  assign v_7636_0 = v_589_0 | v_601_0;
  assign v_7637_0 = v_607_0 | v_26_0;
  assign v_7638_0 = v_7639_0 | v_7977_0;
  assign v_7639_0 = v_7640_0 | v_7976_0;
  assign v_7640_0 = v_589_0 ? v_7641_0 : 3'h0;
  assign v_7642_0 = v_7643_0 | v_7644_0;
  assign v_7643_0 = v_589_0 | v_601_0;
  assign v_7644_0 = v_607_0 | v_26_0;
  assign v_7645_0 = v_7646_0 | v_7973_0;
  assign v_7646_0 = v_7647_0 | v_7972_0;
  assign v_7647_0 = v_589_0 ? v_7648_0 : 3'h0;
  assign v_7649_0 = v_7650_0 | v_7651_0;
  assign v_7650_0 = v_589_0 | v_601_0;
  assign v_7651_0 = v_607_0 | v_26_0;
  assign v_7652_0 = v_7653_0 | v_7969_0;
  assign v_7653_0 = v_7654_0 | v_7968_0;
  assign v_7654_0 = v_589_0 ? v_7655_0 : 3'h0;
  assign v_7656_0 = v_7657_0 | v_7658_0;
  assign v_7657_0 = v_589_0 | v_601_0;
  assign v_7658_0 = v_607_0 | v_26_0;
  assign v_7659_0 = v_7660_0 | v_7965_0;
  assign v_7660_0 = v_7661_0 | v_7964_0;
  assign v_7661_0 = v_589_0 ? v_7662_0 : 3'h0;
  assign v_7663_0 = v_7664_0 | v_7665_0;
  assign v_7664_0 = v_589_0 | v_601_0;
  assign v_7665_0 = v_607_0 | v_26_0;
  assign v_7666_0 = v_7667_0 | v_7961_0;
  assign v_7667_0 = v_7668_0 | v_7960_0;
  assign v_7668_0 = v_589_0 ? v_7669_0 : 3'h0;
  assign v_7670_0 = v_7671_0 | v_7672_0;
  assign v_7671_0 = v_589_0 | v_601_0;
  assign v_7672_0 = v_607_0 | v_26_0;
  assign v_7673_0 = v_7674_0 | v_7957_0;
  assign v_7674_0 = v_7675_0 | v_7956_0;
  assign v_7675_0 = v_589_0 ? v_7676_0 : 3'h0;
  assign v_7677_0 = v_7678_0 | v_7679_0;
  assign v_7678_0 = v_589_0 | v_601_0;
  assign v_7679_0 = v_607_0 | v_26_0;
  assign v_7680_0 = v_7681_0 | v_7953_0;
  assign v_7681_0 = v_7682_0 | v_7952_0;
  assign v_7682_0 = v_589_0 ? v_7683_0 : 3'h0;
  assign v_7684_0 = v_7685_0 | v_7686_0;
  assign v_7685_0 = v_589_0 | v_601_0;
  assign v_7686_0 = v_607_0 | v_26_0;
  assign v_7687_0 = v_7688_0 | v_7949_0;
  assign v_7688_0 = v_7689_0 | v_7948_0;
  assign v_7689_0 = v_589_0 ? v_7690_0 : 3'h0;
  assign v_7691_0 = v_7692_0 | v_7693_0;
  assign v_7692_0 = v_589_0 | v_601_0;
  assign v_7693_0 = v_607_0 | v_26_0;
  assign v_7694_0 = v_7695_0 | v_7945_0;
  assign v_7695_0 = v_7696_0 | v_7944_0;
  assign v_7696_0 = v_589_0 ? v_7697_0 : 3'h0;
  assign v_7698_0 = v_7699_0 | v_7700_0;
  assign v_7699_0 = v_589_0 | v_601_0;
  assign v_7700_0 = v_607_0 | v_26_0;
  assign v_7701_0 = v_7702_0 | v_7941_0;
  assign v_7702_0 = v_7703_0 | v_7940_0;
  assign v_7703_0 = v_589_0 ? v_7704_0 : 3'h0;
  assign v_7705_0 = v_7706_0 | v_7707_0;
  assign v_7706_0 = v_589_0 | v_601_0;
  assign v_7707_0 = v_607_0 | v_26_0;
  assign v_7708_0 = v_7709_0 | v_7937_0;
  assign v_7709_0 = v_7710_0 | v_7936_0;
  assign v_7710_0 = v_589_0 ? v_7711_0 : 3'h0;
  assign v_7712_0 = v_7713_0 | v_7714_0;
  assign v_7713_0 = v_589_0 | v_601_0;
  assign v_7714_0 = v_607_0 | v_26_0;
  assign v_7715_0 = v_7716_0 | v_7933_0;
  assign v_7716_0 = v_7717_0 | v_7932_0;
  assign v_7717_0 = v_589_0 ? v_7718_0 : 3'h0;
  assign v_7719_0 = v_7720_0 | v_7721_0;
  assign v_7720_0 = v_589_0 | v_601_0;
  assign v_7721_0 = v_607_0 | v_26_0;
  assign v_7722_0 = v_7723_0 | v_7929_0;
  assign v_7723_0 = v_7724_0 | v_7928_0;
  assign v_7724_0 = v_589_0 ? v_7725_0 : 3'h0;
  assign v_7726_0 = v_7727_0 | v_7728_0;
  assign v_7727_0 = v_589_0 | v_601_0;
  assign v_7728_0 = v_607_0 | v_26_0;
  assign v_7729_0 = v_7730_0 | v_7925_0;
  assign v_7730_0 = v_7731_0 | v_7924_0;
  assign v_7731_0 = v_589_0 ? v_7732_0 : 3'h0;
  assign v_7733_0 = v_7734_0 | v_7735_0;
  assign v_7734_0 = v_589_0 | v_601_0;
  assign v_7735_0 = v_607_0 | v_26_0;
  assign v_7736_0 = v_7737_0 | v_7921_0;
  assign v_7737_0 = v_7738_0 | v_7920_0;
  assign v_7738_0 = v_589_0 ? v_7739_0 : 3'h0;
  assign v_7740_0 = v_7741_0 | v_7742_0;
  assign v_7741_0 = v_589_0 | v_601_0;
  assign v_7742_0 = v_607_0 | v_26_0;
  assign v_7743_0 = v_7744_0 | v_7917_0;
  assign v_7744_0 = v_7745_0 | v_7916_0;
  assign v_7745_0 = v_589_0 ? v_7746_0 : 3'h0;
  assign v_7747_0 = v_7748_0 | v_7749_0;
  assign v_7748_0 = v_589_0 | v_601_0;
  assign v_7749_0 = v_607_0 | v_26_0;
  assign v_7750_0 = v_7751_0 | v_7913_0;
  assign v_7751_0 = v_7752_0 | v_7912_0;
  assign v_7752_0 = v_589_0 ? v_7753_0 : 3'h0;
  assign v_7754_0 = v_7755_0 | v_7756_0;
  assign v_7755_0 = v_589_0 | v_601_0;
  assign v_7756_0 = v_607_0 | v_26_0;
  assign v_7757_0 = v_7758_0 | v_7909_0;
  assign v_7758_0 = v_7759_0 | v_7908_0;
  assign v_7759_0 = v_589_0 ? v_7760_0 : 3'h0;
  assign v_7761_0 = v_7762_0 | v_7763_0;
  assign v_7762_0 = v_589_0 | v_601_0;
  assign v_7763_0 = v_607_0 | v_26_0;
  assign v_7764_0 = v_7765_0 | v_7905_0;
  assign v_7765_0 = v_7766_0 | v_7904_0;
  assign v_7766_0 = v_589_0 ? v_7767_0 : 3'h0;
  assign v_7768_0 = v_7769_0 | v_7770_0;
  assign v_7769_0 = v_589_0 | v_601_0;
  assign v_7770_0 = v_607_0 | v_26_0;
  assign v_7771_0 = v_7772_0 | v_7901_0;
  assign v_7772_0 = v_7773_0 | v_7900_0;
  assign v_7773_0 = v_589_0 ? v_7774_0 : 3'h0;
  assign v_7775_0 = v_7776_0 | v_7777_0;
  assign v_7776_0 = v_589_0 | v_601_0;
  assign v_7777_0 = v_607_0 | v_26_0;
  assign v_7778_0 = v_7779_0 | v_7897_0;
  assign v_7779_0 = v_7780_0 | v_7896_0;
  assign v_7780_0 = v_589_0 ? v_7781_0 : 3'h0;
  assign v_7782_0 = v_7783_0 | v_7784_0;
  assign v_7783_0 = v_589_0 | v_601_0;
  assign v_7784_0 = v_607_0 | v_26_0;
  assign v_7785_0 = v_7786_0 | v_7893_0;
  assign v_7786_0 = v_7787_0 | v_7892_0;
  assign v_7787_0 = v_589_0 ? v_7788_0 : 3'h0;
  assign v_7789_0 = v_7790_0 | v_7791_0;
  assign v_7790_0 = v_589_0 | v_601_0;
  assign v_7791_0 = v_607_0 | v_26_0;
  assign v_7792_0 = v_7793_0 | v_7889_0;
  assign v_7793_0 = v_7794_0 | v_7888_0;
  assign v_7794_0 = v_589_0 ? v_7795_0 : 3'h0;
  assign v_7796_0 = v_7797_0 | v_7798_0;
  assign v_7797_0 = v_589_0 | v_601_0;
  assign v_7798_0 = v_607_0 | v_26_0;
  assign v_7799_0 = v_7800_0 | v_7885_0;
  assign v_7800_0 = v_7801_0 | v_7884_0;
  assign v_7801_0 = v_589_0 ? v_7802_0 : 3'h0;
  assign v_7803_0 = v_7804_0 | v_7805_0;
  assign v_7804_0 = v_589_0 | v_601_0;
  assign v_7805_0 = v_607_0 | v_26_0;
  assign v_7806_0 = v_7807_0 | v_7881_0;
  assign v_7807_0 = v_7808_0 | v_7880_0;
  assign v_7808_0 = v_589_0 ? v_7809_0 : 3'h0;
  assign v_7810_0 = v_7811_0 | v_7812_0;
  assign v_7811_0 = v_589_0 | v_601_0;
  assign v_7812_0 = v_607_0 | v_26_0;
  assign v_7813_0 = v_7814_0 | v_7877_0;
  assign v_7814_0 = v_7815_0 | v_7876_0;
  assign v_7815_0 = v_589_0 ? v_7816_0 : 3'h0;
  assign v_7817_0 = v_7818_0 | v_7819_0;
  assign v_7818_0 = v_589_0 | v_601_0;
  assign v_7819_0 = v_607_0 | v_26_0;
  assign v_7820_0 = v_7821_0 | v_7873_0;
  assign v_7821_0 = v_7822_0 | v_7872_0;
  assign v_7822_0 = v_589_0 ? v_7823_0 : 3'h0;
  assign v_7824_0 = v_7825_0 | v_7826_0;
  assign v_7825_0 = v_589_0 | v_601_0;
  assign v_7826_0 = v_607_0 | v_26_0;
  assign v_7827_0 = v_7828_0 | v_7869_0;
  assign v_7828_0 = v_7829_0 | v_7868_0;
  assign v_7829_0 = v_589_0 ? v_7830_0 : 3'h0;
  assign v_7831_0 = v_7832_0 | v_7833_0;
  assign v_7832_0 = v_589_0 | v_601_0;
  assign v_7833_0 = v_607_0 | v_26_0;
  assign v_7834_0 = v_7835_0 | v_7865_0;
  assign v_7835_0 = v_7836_0 | v_7864_0;
  assign v_7836_0 = v_589_0 ? v_7837_0 : 3'h0;
  assign v_7838_0 = v_7839_0 | v_7840_0;
  assign v_7839_0 = v_589_0 | v_601_0;
  assign v_7840_0 = v_607_0 | v_26_0;
  assign v_7841_0 = v_7842_0 | v_7861_0;
  assign v_7842_0 = v_7843_0 | v_7860_0;
  assign v_7843_0 = v_589_0 ? v_7844_0 : 3'h0;
  assign v_7845_0 = v_7846_0 | v_7847_0;
  assign v_7846_0 = v_589_0 | v_601_0;
  assign v_7847_0 = v_607_0 | v_26_0;
  assign v_7848_0 = v_7849_0 | v_7857_0;
  assign v_7849_0 = v_7850_0 | v_7856_0;
  assign v_7850_0 = v_589_0 ? v_7851_0 : 3'h0;
  assign v_7852_0 = v_601_0 | v_26_0;
  assign v_7853_0 = v_7854_0 | v_7855_0;
  assign v_7854_0 = v_601_0 ? v_7844_0 : 3'h0;
  assign v_7855_0 = v_26_0 ? v_7844_0 : 3'h0;
  assign v_7856_0 = v_601_0 ? v_7837_0 : 3'h0;
  assign v_7857_0 = v_7858_0 | v_7859_0;
  assign v_7858_0 = v_607_0 ? v_7851_0 : 3'h0;
  assign v_7859_0 = v_26_0 ? v_7837_0 : 3'h0;
  assign v_7860_0 = v_601_0 ? v_7830_0 : 3'h0;
  assign v_7861_0 = v_7862_0 | v_7863_0;
  assign v_7862_0 = v_607_0 ? v_7844_0 : 3'h0;
  assign v_7863_0 = v_26_0 ? v_7830_0 : 3'h0;
  assign v_7864_0 = v_601_0 ? v_7823_0 : 3'h0;
  assign v_7865_0 = v_7866_0 | v_7867_0;
  assign v_7866_0 = v_607_0 ? v_7837_0 : 3'h0;
  assign v_7867_0 = v_26_0 ? v_7823_0 : 3'h0;
  assign v_7868_0 = v_601_0 ? v_7816_0 : 3'h0;
  assign v_7869_0 = v_7870_0 | v_7871_0;
  assign v_7870_0 = v_607_0 ? v_7830_0 : 3'h0;
  assign v_7871_0 = v_26_0 ? v_7816_0 : 3'h0;
  assign v_7872_0 = v_601_0 ? v_7809_0 : 3'h0;
  assign v_7873_0 = v_7874_0 | v_7875_0;
  assign v_7874_0 = v_607_0 ? v_7823_0 : 3'h0;
  assign v_7875_0 = v_26_0 ? v_7809_0 : 3'h0;
  assign v_7876_0 = v_601_0 ? v_7802_0 : 3'h0;
  assign v_7877_0 = v_7878_0 | v_7879_0;
  assign v_7878_0 = v_607_0 ? v_7816_0 : 3'h0;
  assign v_7879_0 = v_26_0 ? v_7802_0 : 3'h0;
  assign v_7880_0 = v_601_0 ? v_7795_0 : 3'h0;
  assign v_7881_0 = v_7882_0 | v_7883_0;
  assign v_7882_0 = v_607_0 ? v_7809_0 : 3'h0;
  assign v_7883_0 = v_26_0 ? v_7795_0 : 3'h0;
  assign v_7884_0 = v_601_0 ? v_7788_0 : 3'h0;
  assign v_7885_0 = v_7886_0 | v_7887_0;
  assign v_7886_0 = v_607_0 ? v_7802_0 : 3'h0;
  assign v_7887_0 = v_26_0 ? v_7788_0 : 3'h0;
  assign v_7888_0 = v_601_0 ? v_7781_0 : 3'h0;
  assign v_7889_0 = v_7890_0 | v_7891_0;
  assign v_7890_0 = v_607_0 ? v_7795_0 : 3'h0;
  assign v_7891_0 = v_26_0 ? v_7781_0 : 3'h0;
  assign v_7892_0 = v_601_0 ? v_7774_0 : 3'h0;
  assign v_7893_0 = v_7894_0 | v_7895_0;
  assign v_7894_0 = v_607_0 ? v_7788_0 : 3'h0;
  assign v_7895_0 = v_26_0 ? v_7774_0 : 3'h0;
  assign v_7896_0 = v_601_0 ? v_7767_0 : 3'h0;
  assign v_7897_0 = v_7898_0 | v_7899_0;
  assign v_7898_0 = v_607_0 ? v_7781_0 : 3'h0;
  assign v_7899_0 = v_26_0 ? v_7767_0 : 3'h0;
  assign v_7900_0 = v_601_0 ? v_7760_0 : 3'h0;
  assign v_7901_0 = v_7902_0 | v_7903_0;
  assign v_7902_0 = v_607_0 ? v_7774_0 : 3'h0;
  assign v_7903_0 = v_26_0 ? v_7760_0 : 3'h0;
  assign v_7904_0 = v_601_0 ? v_7753_0 : 3'h0;
  assign v_7905_0 = v_7906_0 | v_7907_0;
  assign v_7906_0 = v_607_0 ? v_7767_0 : 3'h0;
  assign v_7907_0 = v_26_0 ? v_7753_0 : 3'h0;
  assign v_7908_0 = v_601_0 ? v_7746_0 : 3'h0;
  assign v_7909_0 = v_7910_0 | v_7911_0;
  assign v_7910_0 = v_607_0 ? v_7760_0 : 3'h0;
  assign v_7911_0 = v_26_0 ? v_7746_0 : 3'h0;
  assign v_7912_0 = v_601_0 ? v_7739_0 : 3'h0;
  assign v_7913_0 = v_7914_0 | v_7915_0;
  assign v_7914_0 = v_607_0 ? v_7753_0 : 3'h0;
  assign v_7915_0 = v_26_0 ? v_7739_0 : 3'h0;
  assign v_7916_0 = v_601_0 ? v_7732_0 : 3'h0;
  assign v_7917_0 = v_7918_0 | v_7919_0;
  assign v_7918_0 = v_607_0 ? v_7746_0 : 3'h0;
  assign v_7919_0 = v_26_0 ? v_7732_0 : 3'h0;
  assign v_7920_0 = v_601_0 ? v_7725_0 : 3'h0;
  assign v_7921_0 = v_7922_0 | v_7923_0;
  assign v_7922_0 = v_607_0 ? v_7739_0 : 3'h0;
  assign v_7923_0 = v_26_0 ? v_7725_0 : 3'h0;
  assign v_7924_0 = v_601_0 ? v_7718_0 : 3'h0;
  assign v_7925_0 = v_7926_0 | v_7927_0;
  assign v_7926_0 = v_607_0 ? v_7732_0 : 3'h0;
  assign v_7927_0 = v_26_0 ? v_7718_0 : 3'h0;
  assign v_7928_0 = v_601_0 ? v_7711_0 : 3'h0;
  assign v_7929_0 = v_7930_0 | v_7931_0;
  assign v_7930_0 = v_607_0 ? v_7725_0 : 3'h0;
  assign v_7931_0 = v_26_0 ? v_7711_0 : 3'h0;
  assign v_7932_0 = v_601_0 ? v_7704_0 : 3'h0;
  assign v_7933_0 = v_7934_0 | v_7935_0;
  assign v_7934_0 = v_607_0 ? v_7718_0 : 3'h0;
  assign v_7935_0 = v_26_0 ? v_7704_0 : 3'h0;
  assign v_7936_0 = v_601_0 ? v_7697_0 : 3'h0;
  assign v_7937_0 = v_7938_0 | v_7939_0;
  assign v_7938_0 = v_607_0 ? v_7711_0 : 3'h0;
  assign v_7939_0 = v_26_0 ? v_7697_0 : 3'h0;
  assign v_7940_0 = v_601_0 ? v_7690_0 : 3'h0;
  assign v_7941_0 = v_7942_0 | v_7943_0;
  assign v_7942_0 = v_607_0 ? v_7704_0 : 3'h0;
  assign v_7943_0 = v_26_0 ? v_7690_0 : 3'h0;
  assign v_7944_0 = v_601_0 ? v_7683_0 : 3'h0;
  assign v_7945_0 = v_7946_0 | v_7947_0;
  assign v_7946_0 = v_607_0 ? v_7697_0 : 3'h0;
  assign v_7947_0 = v_26_0 ? v_7683_0 : 3'h0;
  assign v_7948_0 = v_601_0 ? v_7676_0 : 3'h0;
  assign v_7949_0 = v_7950_0 | v_7951_0;
  assign v_7950_0 = v_607_0 ? v_7690_0 : 3'h0;
  assign v_7951_0 = v_26_0 ? v_7676_0 : 3'h0;
  assign v_7952_0 = v_601_0 ? v_7669_0 : 3'h0;
  assign v_7953_0 = v_7954_0 | v_7955_0;
  assign v_7954_0 = v_607_0 ? v_7683_0 : 3'h0;
  assign v_7955_0 = v_26_0 ? v_7669_0 : 3'h0;
  assign v_7956_0 = v_601_0 ? v_7662_0 : 3'h0;
  assign v_7957_0 = v_7958_0 | v_7959_0;
  assign v_7958_0 = v_607_0 ? v_7676_0 : 3'h0;
  assign v_7959_0 = v_26_0 ? v_7662_0 : 3'h0;
  assign v_7960_0 = v_601_0 ? v_7655_0 : 3'h0;
  assign v_7961_0 = v_7962_0 | v_7963_0;
  assign v_7962_0 = v_607_0 ? v_7669_0 : 3'h0;
  assign v_7963_0 = v_26_0 ? v_7655_0 : 3'h0;
  assign v_7964_0 = v_601_0 ? v_7648_0 : 3'h0;
  assign v_7965_0 = v_7966_0 | v_7967_0;
  assign v_7966_0 = v_607_0 ? v_7662_0 : 3'h0;
  assign v_7967_0 = v_26_0 ? v_7648_0 : 3'h0;
  assign v_7968_0 = v_601_0 ? v_7641_0 : 3'h0;
  assign v_7969_0 = v_7970_0 | v_7971_0;
  assign v_7970_0 = v_607_0 ? v_7655_0 : 3'h0;
  assign v_7971_0 = v_26_0 ? v_7641_0 : 3'h0;
  assign v_7972_0 = v_601_0 ? v_7634_0 : 3'h0;
  assign v_7973_0 = v_7974_0 | v_7975_0;
  assign v_7974_0 = v_607_0 ? v_7648_0 : 3'h0;
  assign v_7975_0 = v_26_0 ? v_7634_0 : 3'h0;
  assign v_7976_0 = v_601_0 ? v_7627_0 : 3'h0;
  assign v_7977_0 = v_7978_0 | v_7979_0;
  assign v_7978_0 = v_607_0 ? v_7641_0 : 3'h0;
  assign v_7979_0 = v_26_0 ? v_7627_0 : 3'h0;
  assign v_7980_0 = v_601_0 ? v_7620_0 : 3'h0;
  assign v_7981_0 = v_7982_0 | v_7983_0;
  assign v_7982_0 = v_607_0 ? v_7634_0 : 3'h0;
  assign v_7983_0 = v_26_0 ? v_7620_0 : 3'h0;
  assign v_7984_0 = v_601_0 ? v_7613_0 : 3'h0;
  assign v_7985_0 = v_7986_0 | v_7987_0;
  assign v_7986_0 = v_607_0 ? v_7627_0 : 3'h0;
  assign v_7987_0 = v_26_0 ? v_7613_0 : 3'h0;
  assign v_7988_0 = v_601_0 ? v_7606_0 : 3'h0;
  assign v_7989_0 = v_7990_0 | v_7991_0;
  assign v_7990_0 = v_607_0 ? v_7620_0 : 3'h0;
  assign v_7991_0 = v_26_0 ? v_7606_0 : 3'h0;
  assign v_7992_0 = v_601_0 ? v_7599_0 : 3'h0;
  assign v_7993_0 = v_7994_0 | v_7995_0;
  assign v_7994_0 = v_607_0 ? v_7613_0 : 3'h0;
  assign v_7995_0 = v_26_0 ? v_7599_0 : 3'h0;
  assign v_7996_0 = v_601_0 ? v_7592_0 : 3'h0;
  assign v_7997_0 = v_7998_0 | v_7999_0;
  assign v_7998_0 = v_607_0 ? v_7606_0 : 3'h0;
  assign v_7999_0 = v_26_0 ? v_7592_0 : 3'h0;
  assign v_8000_0 = v_601_0 ? v_7585_0 : 3'h0;
  assign v_8001_0 = v_8002_0 | v_8003_0;
  assign v_8002_0 = v_607_0 ? v_7599_0 : 3'h0;
  assign v_8003_0 = v_26_0 ? v_7585_0 : 3'h0;
  assign v_8004_0 = v_601_0 ? v_7578_0 : 3'h0;
  assign v_8005_0 = v_8006_0 | v_8007_0;
  assign v_8006_0 = v_607_0 ? v_7592_0 : 3'h0;
  assign v_8007_0 = v_26_0 ? v_7578_0 : 3'h0;
  assign v_8008_0 = v_601_0 ? v_7571_0 : 3'h0;
  assign v_8009_0 = v_8010_0 | v_8011_0;
  assign v_8010_0 = v_607_0 ? v_7585_0 : 3'h0;
  assign v_8011_0 = v_26_0 ? v_7571_0 : 3'h0;
  assign v_8012_0 = v_601_0 ? v_7564_0 : 3'h0;
  assign v_8013_0 = v_8014_0 | v_8015_0;
  assign v_8014_0 = v_607_0 ? v_7578_0 : 3'h0;
  assign v_8015_0 = v_26_0 ? v_7564_0 : 3'h0;
  assign v_8016_0 = v_601_0 ? v_7557_0 : 3'h0;
  assign v_8017_0 = v_8018_0 | v_8019_0;
  assign v_8018_0 = v_607_0 ? v_7571_0 : 3'h0;
  assign v_8019_0 = v_26_0 ? v_7557_0 : 3'h0;
  assign v_8020_0 = v_601_0 ? v_7550_0 : 3'h0;
  assign v_8021_0 = v_8022_0 | v_8023_0;
  assign v_8022_0 = v_607_0 ? v_7564_0 : 3'h0;
  assign v_8023_0 = v_26_0 ? v_7550_0 : 3'h0;
  assign v_8024_0 = v_601_0 ? v_7543_0 : 3'h0;
  assign v_8025_0 = v_8026_0 | v_8027_0;
  assign v_8026_0 = v_607_0 ? v_7557_0 : 3'h0;
  assign v_8027_0 = v_26_0 ? v_7543_0 : 3'h0;
  assign v_8028_0 = v_601_0 ? v_7536_0 : 3'h0;
  assign v_8029_0 = v_8030_0 | v_8031_0;
  assign v_8030_0 = v_607_0 ? v_7550_0 : 3'h0;
  assign v_8031_0 = v_26_0 ? v_7536_0 : 3'h0;
  assign v_8032_0 = v_601_0 ? v_7529_0 : 3'h0;
  assign v_8033_0 = v_8034_0 | v_8035_0;
  assign v_8034_0 = v_607_0 ? v_7543_0 : 3'h0;
  assign v_8035_0 = v_26_0 ? v_7529_0 : 3'h0;
  assign v_8036_0 = v_601_0 ? v_7522_0 : 3'h0;
  assign v_8037_0 = v_8038_0 | v_8039_0;
  assign v_8038_0 = v_607_0 ? v_7536_0 : 3'h0;
  assign v_8039_0 = v_26_0 ? v_7522_0 : 3'h0;
  assign v_8040_0 = v_601_0 ? v_7515_0 : 3'h0;
  assign v_8041_0 = v_8042_0 | v_8043_0;
  assign v_8042_0 = v_607_0 ? v_7529_0 : 3'h0;
  assign v_8043_0 = v_26_0 ? v_7515_0 : 3'h0;
  assign v_8044_0 = v_601_0 ? v_7508_0 : 3'h0;
  assign v_8045_0 = v_8046_0 | v_8047_0;
  assign v_8046_0 = v_607_0 ? v_7522_0 : 3'h0;
  assign v_8047_0 = v_26_0 ? v_7508_0 : 3'h0;
  assign v_8048_0 = v_601_0 ? v_7501_0 : 3'h0;
  assign v_8049_0 = v_8050_0 | v_8051_0;
  assign v_8050_0 = v_607_0 ? v_7515_0 : 3'h0;
  assign v_8051_0 = v_26_0 ? v_7501_0 : 3'h0;
  assign v_8052_0 = v_601_0 ? v_7494_0 : 3'h0;
  assign v_8053_0 = v_8054_0 | v_8055_0;
  assign v_8054_0 = v_607_0 ? v_7508_0 : 3'h0;
  assign v_8055_0 = v_26_0 ? v_7494_0 : 3'h0;
  assign v_8056_0 = v_601_0 ? v_7487_0 : 3'h0;
  assign v_8057_0 = v_8058_0 | v_8059_0;
  assign v_8058_0 = v_607_0 ? v_7501_0 : 3'h0;
  assign v_8059_0 = v_26_0 ? v_7487_0 : 3'h0;
  assign v_8060_0 = v_601_0 ? v_7480_0 : 3'h0;
  assign v_8061_0 = v_8062_0 | v_8063_0;
  assign v_8062_0 = v_607_0 ? v_7494_0 : 3'h0;
  assign v_8063_0 = v_26_0 ? v_7480_0 : 3'h0;
  assign v_8064_0 = v_601_0 ? v_7473_0 : 3'h0;
  assign v_8065_0 = v_8066_0 | v_8067_0;
  assign v_8066_0 = v_607_0 ? v_7487_0 : 3'h0;
  assign v_8067_0 = v_26_0 ? v_7473_0 : 3'h0;
  assign v_8068_0 = v_601_0 ? v_7466_0 : 3'h0;
  assign v_8069_0 = v_8070_0 | v_8071_0;
  assign v_8070_0 = v_607_0 ? v_7480_0 : 3'h0;
  assign v_8071_0 = v_26_0 ? v_7466_0 : 3'h0;
  assign v_8072_0 = v_601_0 ? v_7459_0 : 3'h0;
  assign v_8073_0 = v_8074_0 | v_8075_0;
  assign v_8074_0 = v_607_0 ? v_7473_0 : 3'h0;
  assign v_8075_0 = v_26_0 ? v_7459_0 : 3'h0;
  assign v_8076_0 = v_601_0 ? v_7452_0 : 3'h0;
  assign v_8077_0 = v_8078_0 | v_8079_0;
  assign v_8078_0 = v_607_0 ? v_7466_0 : 3'h0;
  assign v_8079_0 = v_26_0 ? v_7452_0 : 3'h0;
  assign v_8080_0 = v_601_0 ? v_7445_0 : 3'h0;
  assign v_8081_0 = v_8082_0 | v_8083_0;
  assign v_8082_0 = v_607_0 ? v_7459_0 : 3'h0;
  assign v_8083_0 = v_26_0 ? v_7445_0 : 3'h0;
  assign v_8084_0 = v_601_0 ? v_7438_0 : 3'h0;
  assign v_8085_0 = v_8086_0 | v_8087_0;
  assign v_8086_0 = v_607_0 ? v_7452_0 : 3'h0;
  assign v_8087_0 = v_26_0 ? v_7438_0 : 3'h0;
  assign v_8088_0 = v_601_0 ? v_7431_0 : 3'h0;
  assign v_8089_0 = v_8090_0 | v_8091_0;
  assign v_8090_0 = v_607_0 ? v_7445_0 : 3'h0;
  assign v_8091_0 = v_26_0 ? v_7431_0 : 3'h0;
  assign v_8092_0 = v_601_0 ? v_7424_0 : 3'h0;
  assign v_8093_0 = v_8094_0 | v_8095_0;
  assign v_8094_0 = v_607_0 ? v_7438_0 : 3'h0;
  assign v_8095_0 = v_26_0 ? v_7424_0 : 3'h0;
  assign v_8096_0 = v_601_0 ? v_7417_0 : 3'h0;
  assign v_8097_0 = v_8098_0 | v_8099_0;
  assign v_8098_0 = v_607_0 ? v_7431_0 : 3'h0;
  assign v_8099_0 = v_26_0 ? v_7417_0 : 3'h0;
  assign v_8100_0 = v_601_0 ? v_7410_0 : 3'h0;
  assign v_8101_0 = v_8102_0 | v_8103_0;
  assign v_8102_0 = v_607_0 ? v_7424_0 : 3'h0;
  assign v_8103_0 = v_26_0 ? v_7410_0 : 3'h0;
  assign v_8104_0 = v_601_0 ? v_7403_0 : 3'h0;
  assign v_8105_0 = v_8106_0 | v_8107_0;
  assign v_8106_0 = v_607_0 ? v_7417_0 : 3'h0;
  assign v_8107_0 = v_26_0 ? v_7403_0 : 3'h0;
  assign v_8108_0 = v_601_0 ? v_7396_0 : 3'h0;
  assign v_8109_0 = v_8110_0 | v_8111_0;
  assign v_8110_0 = v_607_0 ? v_7410_0 : 3'h0;
  assign v_8111_0 = v_26_0 ? v_7396_0 : 3'h0;
  assign v_8112_0 = v_601_0 ? v_7389_0 : 3'h0;
  assign v_8113_0 = v_8114_0 | v_8115_0;
  assign v_8114_0 = v_607_0 ? v_7403_0 : 3'h0;
  assign v_8115_0 = v_26_0 ? v_7389_0 : 3'h0;
  assign v_8116_0 = v_601_0 ? v_7382_0 : 3'h0;
  assign v_8117_0 = v_8118_0 | v_8119_0;
  assign v_8118_0 = v_607_0 ? v_7396_0 : 3'h0;
  assign v_8119_0 = v_26_0 ? v_7382_0 : 3'h0;
  assign v_8120_0 = v_601_0 ? v_7375_0 : 3'h0;
  assign v_8121_0 = v_8122_0 | v_8123_0;
  assign v_8122_0 = v_607_0 ? v_7389_0 : 3'h0;
  assign v_8123_0 = v_26_0 ? v_7375_0 : 3'h0;
  assign v_8124_0 = v_601_0 ? v_7368_0 : 3'h0;
  assign v_8125_0 = v_8126_0 | v_8127_0;
  assign v_8126_0 = v_607_0 ? v_7382_0 : 3'h0;
  assign v_8127_0 = v_26_0 ? v_7368_0 : 3'h0;
  assign v_8128_0 = v_601_0 ? v_7361_0 : 3'h0;
  assign v_8129_0 = v_8130_0 | v_8131_0;
  assign v_8130_0 = v_607_0 ? v_7375_0 : 3'h0;
  assign v_8131_0 = v_26_0 ? v_7361_0 : 3'h0;
  assign v_8132_0 = v_601_0 ? v_7354_0 : 3'h0;
  assign v_8133_0 = v_8134_0 | v_8135_0;
  assign v_8134_0 = v_607_0 ? v_7368_0 : 3'h0;
  assign v_8135_0 = v_26_0 ? v_7354_0 : 3'h0;
  assign v_8136_0 = v_601_0 ? v_7347_0 : 3'h0;
  assign v_8137_0 = v_8138_0 | v_8139_0;
  assign v_8138_0 = v_607_0 ? v_7361_0 : 3'h0;
  assign v_8139_0 = v_26_0 ? v_7347_0 : 3'h0;
  assign v_8140_0 = v_601_0 ? v_7340_0 : 3'h0;
  assign v_8141_0 = v_8142_0 | v_8143_0;
  assign v_8142_0 = v_607_0 ? v_7354_0 : 3'h0;
  assign v_8143_0 = v_26_0 ? v_7340_0 : 3'h0;
  assign v_8144_0 = v_601_0 ? v_7333_0 : 3'h0;
  assign v_8145_0 = v_8146_0 | v_8147_0;
  assign v_8146_0 = v_607_0 ? v_7347_0 : 3'h0;
  assign v_8147_0 = v_26_0 ? v_7333_0 : 3'h0;
  assign v_8148_0 = v_601_0 ? v_7326_0 : 3'h0;
  assign v_8149_0 = v_8150_0 | v_8151_0;
  assign v_8150_0 = v_607_0 ? v_7340_0 : 3'h0;
  assign v_8151_0 = v_26_0 ? v_7326_0 : 3'h0;
  assign v_8152_0 = v_601_0 ? v_7319_0 : 3'h0;
  assign v_8153_0 = v_8154_0 | v_8155_0;
  assign v_8154_0 = v_607_0 ? v_7333_0 : 3'h0;
  assign v_8155_0 = v_26_0 ? v_7319_0 : 3'h0;
  assign v_8156_0 = v_601_0 ? v_7312_0 : 3'h0;
  assign v_8157_0 = v_8158_0 | v_8159_0;
  assign v_8158_0 = v_607_0 ? v_7326_0 : 3'h0;
  assign v_8159_0 = v_26_0 ? v_7312_0 : 3'h0;
  assign v_8160_0 = v_601_0 ? v_7305_0 : 3'h0;
  assign v_8161_0 = v_8162_0 | v_8163_0;
  assign v_8162_0 = v_607_0 ? v_7319_0 : 3'h0;
  assign v_8163_0 = v_26_0 ? v_7305_0 : 3'h0;
  assign v_8164_0 = v_601_0 ? v_7298_0 : 3'h0;
  assign v_8165_0 = v_8166_0 | v_8167_0;
  assign v_8166_0 = v_607_0 ? v_7312_0 : 3'h0;
  assign v_8167_0 = v_26_0 ? v_7298_0 : 3'h0;
  assign v_8168_0 = v_601_0 ? v_7291_0 : 3'h0;
  assign v_8169_0 = v_8170_0 | v_8171_0;
  assign v_8170_0 = v_607_0 ? v_7305_0 : 3'h0;
  assign v_8171_0 = v_26_0 ? v_7291_0 : 3'h0;
  assign v_8172_0 = v_601_0 ? v_7284_0 : 3'h0;
  assign v_8173_0 = v_8174_0 | v_8175_0;
  assign v_8174_0 = v_607_0 ? v_7298_0 : 3'h0;
  assign v_8175_0 = v_26_0 ? v_7284_0 : 3'h0;
  assign v_8176_0 = v_601_0 ? v_7277_0 : 3'h0;
  assign v_8177_0 = v_8178_0 | v_8179_0;
  assign v_8178_0 = v_607_0 ? v_7291_0 : 3'h0;
  assign v_8179_0 = v_26_0 ? v_7277_0 : 3'h0;
  assign v_8180_0 = v_601_0 ? v_7270_0 : 3'h0;
  assign v_8181_0 = v_8182_0 | v_8183_0;
  assign v_8182_0 = v_607_0 ? v_7284_0 : 3'h0;
  assign v_8183_0 = v_26_0 ? v_7270_0 : 3'h0;
  assign v_8184_0 = v_601_0 ? v_7263_0 : 3'h0;
  assign v_8185_0 = v_8186_0 | v_8187_0;
  assign v_8186_0 = v_607_0 ? v_7277_0 : 3'h0;
  assign v_8187_0 = v_26_0 ? v_7263_0 : 3'h0;
  assign v_8188_0 = v_601_0 ? v_7256_0 : 3'h0;
  assign v_8189_0 = v_8190_0 | v_8191_0;
  assign v_8190_0 = v_607_0 ? v_7270_0 : 3'h0;
  assign v_8191_0 = v_26_0 ? v_7256_0 : 3'h0;
  assign v_8192_0 = v_601_0 ? v_7249_0 : 3'h0;
  assign v_8193_0 = v_8194_0 | v_8195_0;
  assign v_8194_0 = v_607_0 ? v_7263_0 : 3'h0;
  assign v_8195_0 = v_26_0 ? v_7249_0 : 3'h0;
  assign v_8196_0 = v_601_0 ? v_7242_0 : 3'h0;
  assign v_8197_0 = v_8198_0 | v_8199_0;
  assign v_8198_0 = v_607_0 ? v_7256_0 : 3'h0;
  assign v_8199_0 = v_26_0 ? v_7242_0 : 3'h0;
  assign v_8200_0 = v_601_0 ? v_7235_0 : 3'h0;
  assign v_8201_0 = v_8202_0 | v_8203_0;
  assign v_8202_0 = v_607_0 ? v_7249_0 : 3'h0;
  assign v_8203_0 = v_26_0 ? v_7235_0 : 3'h0;
  assign v_8204_0 = v_601_0 ? v_7228_0 : 3'h0;
  assign v_8205_0 = v_8206_0 | v_8207_0;
  assign v_8206_0 = v_607_0 ? v_7242_0 : 3'h0;
  assign v_8207_0 = v_26_0 ? v_7228_0 : 3'h0;
  assign v_8208_0 = v_601_0 ? v_7221_0 : 3'h0;
  assign v_8209_0 = v_8210_0 | v_8211_0;
  assign v_8210_0 = v_607_0 ? v_7235_0 : 3'h0;
  assign v_8211_0 = v_26_0 ? v_7221_0 : 3'h0;
  assign v_8212_0 = v_601_0 ? v_7214_0 : 3'h0;
  assign v_8213_0 = v_8214_0 | v_8215_0;
  assign v_8214_0 = v_607_0 ? v_7228_0 : 3'h0;
  assign v_8215_0 = v_26_0 ? v_7214_0 : 3'h0;
  assign v_8216_0 = v_601_0 ? v_7207_0 : 3'h0;
  assign v_8217_0 = v_8218_0 | v_8219_0;
  assign v_8218_0 = v_607_0 ? v_7221_0 : 3'h0;
  assign v_8219_0 = v_26_0 ? v_7207_0 : 3'h0;
  assign v_8220_0 = v_601_0 ? v_7200_0 : 3'h0;
  assign v_8221_0 = v_8222_0 | v_8223_0;
  assign v_8222_0 = v_607_0 ? v_7214_0 : 3'h0;
  assign v_8223_0 = v_26_0 ? v_7200_0 : 3'h0;
  assign v_8224_0 = v_601_0 ? v_7193_0 : 3'h0;
  assign v_8225_0 = v_8226_0 | v_8227_0;
  assign v_8226_0 = v_607_0 ? v_7207_0 : 3'h0;
  assign v_8227_0 = v_26_0 ? v_7193_0 : 3'h0;
  assign v_8228_0 = v_601_0 ? v_7186_0 : 3'h0;
  assign v_8229_0 = v_8230_0 | v_8231_0;
  assign v_8230_0 = v_607_0 ? v_7200_0 : 3'h0;
  assign v_8231_0 = v_26_0 ? v_7186_0 : 3'h0;
  assign v_8232_0 = v_601_0 ? v_7179_0 : 3'h0;
  assign v_8233_0 = v_8234_0 | v_8235_0;
  assign v_8234_0 = v_607_0 ? v_7193_0 : 3'h0;
  assign v_8235_0 = v_26_0 ? v_7179_0 : 3'h0;
  assign v_8236_0 = v_601_0 ? v_7172_0 : 3'h0;
  assign v_8237_0 = v_8238_0 | v_8239_0;
  assign v_8238_0 = v_607_0 ? v_7186_0 : 3'h0;
  assign v_8239_0 = v_26_0 ? v_7172_0 : 3'h0;
  assign v_8240_0 = v_601_0 ? v_7165_0 : 3'h0;
  assign v_8241_0 = v_8242_0 | v_8243_0;
  assign v_8242_0 = v_607_0 ? v_7179_0 : 3'h0;
  assign v_8243_0 = v_26_0 ? v_7165_0 : 3'h0;
  assign v_8244_0 = v_601_0 ? v_7158_0 : 3'h0;
  assign v_8245_0 = v_8246_0 | v_8247_0;
  assign v_8246_0 = v_607_0 ? v_7172_0 : 3'h0;
  assign v_8247_0 = v_26_0 ? v_7158_0 : 3'h0;
  assign v_8248_0 = v_601_0 ? v_7151_0 : 3'h0;
  assign v_8249_0 = v_8250_0 | v_8251_0;
  assign v_8250_0 = v_607_0 ? v_7165_0 : 3'h0;
  assign v_8251_0 = v_26_0 ? v_7151_0 : 3'h0;
  assign v_8252_0 = v_601_0 ? v_7144_0 : 3'h0;
  assign v_8253_0 = v_8254_0 | v_8255_0;
  assign v_8254_0 = v_607_0 ? v_7158_0 : 3'h0;
  assign v_8255_0 = v_26_0 ? v_7144_0 : 3'h0;
  assign v_8256_0 = v_601_0 ? v_7137_0 : 3'h0;
  assign v_8257_0 = v_8258_0 | v_8259_0;
  assign v_8258_0 = v_607_0 ? v_7151_0 : 3'h0;
  assign v_8259_0 = v_26_0 ? v_7137_0 : 3'h0;
  assign v_8260_0 = v_601_0 ? v_7130_0 : 3'h0;
  assign v_8261_0 = v_8262_0 | v_8263_0;
  assign v_8262_0 = v_607_0 ? v_7144_0 : 3'h0;
  assign v_8263_0 = v_26_0 ? v_7130_0 : 3'h0;
  assign v_8264_0 = v_601_0 ? v_7123_0 : 3'h0;
  assign v_8265_0 = v_8266_0 | v_8267_0;
  assign v_8266_0 = v_607_0 ? v_7137_0 : 3'h0;
  assign v_8267_0 = v_26_0 ? v_7123_0 : 3'h0;
  assign v_8268_0 = v_601_0 ? v_7116_0 : 3'h0;
  assign v_8269_0 = v_8270_0 | v_8271_0;
  assign v_8270_0 = v_607_0 ? v_7130_0 : 3'h0;
  assign v_8271_0 = v_26_0 ? v_7116_0 : 3'h0;
  assign v_8272_0 = v_601_0 ? v_7109_0 : 3'h0;
  assign v_8273_0 = v_8274_0 | v_8275_0;
  assign v_8274_0 = v_607_0 ? v_7123_0 : 3'h0;
  assign v_8275_0 = v_26_0 ? v_7109_0 : 3'h0;
  assign v_8276_0 = v_601_0 ? v_7102_0 : 3'h0;
  assign v_8277_0 = v_8278_0 | v_8279_0;
  assign v_8278_0 = v_607_0 ? v_7116_0 : 3'h0;
  assign v_8279_0 = v_26_0 ? v_7102_0 : 3'h0;
  assign v_8280_0 = v_601_0 ? v_7095_0 : 3'h0;
  assign v_8281_0 = v_8282_0 | v_8283_0;
  assign v_8282_0 = v_607_0 ? v_7109_0 : 3'h0;
  assign v_8283_0 = v_26_0 ? v_7095_0 : 3'h0;
  assign v_8284_0 = v_601_0 ? v_7088_0 : 3'h0;
  assign v_8285_0 = v_8286_0 | v_8287_0;
  assign v_8286_0 = v_607_0 ? v_7102_0 : 3'h0;
  assign v_8287_0 = v_26_0 ? v_7088_0 : 3'h0;
  assign v_8288_0 = v_601_0 ? v_7081_0 : 3'h0;
  assign v_8289_0 = v_8290_0 | v_8291_0;
  assign v_8290_0 = v_607_0 ? v_7095_0 : 3'h0;
  assign v_8291_0 = v_26_0 ? v_7081_0 : 3'h0;
  assign v_8292_0 = v_601_0 ? v_7074_0 : 3'h0;
  assign v_8293_0 = v_8294_0 | v_8295_0;
  assign v_8294_0 = v_607_0 ? v_7088_0 : 3'h0;
  assign v_8295_0 = v_26_0 ? v_7074_0 : 3'h0;
  assign v_8296_0 = v_601_0 ? v_7067_0 : 3'h0;
  assign v_8297_0 = v_8298_0 | v_8299_0;
  assign v_8298_0 = v_607_0 ? v_7081_0 : 3'h0;
  assign v_8299_0 = v_26_0 ? v_7067_0 : 3'h0;
  assign v_8300_0 = v_601_0 ? v_7060_0 : 3'h0;
  assign v_8301_0 = v_8302_0 | v_8303_0;
  assign v_8302_0 = v_607_0 ? v_7074_0 : 3'h0;
  assign v_8303_0 = v_26_0 ? v_7060_0 : 3'h0;
  assign v_8304_0 = v_601_0 ? v_7053_0 : 3'h0;
  assign v_8305_0 = v_8306_0 | v_8307_0;
  assign v_8306_0 = v_607_0 ? v_7067_0 : 3'h0;
  assign v_8307_0 = v_26_0 ? v_7053_0 : 3'h0;
  assign v_8308_0 = v_601_0 ? v_7046_0 : 3'h0;
  assign v_8309_0 = v_8310_0 | v_8311_0;
  assign v_8310_0 = v_607_0 ? v_7060_0 : 3'h0;
  assign v_8311_0 = v_26_0 ? v_7046_0 : 3'h0;
  assign v_8312_0 = v_601_0 ? v_7039_0 : 3'h0;
  assign v_8313_0 = v_8314_0 | v_8315_0;
  assign v_8314_0 = v_607_0 ? v_7053_0 : 3'h0;
  assign v_8315_0 = v_26_0 ? v_7039_0 : 3'h0;
  assign v_8316_0 = v_601_0 ? v_7032_0 : 3'h0;
  assign v_8317_0 = v_8318_0 | v_8319_0;
  assign v_8318_0 = v_607_0 ? v_7046_0 : 3'h0;
  assign v_8319_0 = v_26_0 ? v_7032_0 : 3'h0;
  assign v_8320_0 = v_601_0 ? v_7025_0 : 3'h0;
  assign v_8321_0 = v_8322_0 | v_8323_0;
  assign v_8322_0 = v_607_0 ? v_7039_0 : 3'h0;
  assign v_8323_0 = v_26_0 ? v_7025_0 : 3'h0;
  assign v_8324_0 = v_601_0 ? v_7018_0 : 3'h0;
  assign v_8325_0 = v_8326_0 | v_8327_0;
  assign v_8326_0 = v_607_0 ? v_7032_0 : 3'h0;
  assign v_8327_0 = v_26_0 ? v_7018_0 : 3'h0;
  assign v_8328_0 = v_601_0 ? v_7011_0 : 3'h0;
  assign v_8329_0 = v_8330_0 | v_8331_0;
  assign v_8330_0 = v_607_0 ? v_7025_0 : 3'h0;
  assign v_8331_0 = v_26_0 ? v_7011_0 : 3'h0;
  assign v_8332_0 = v_601_0 ? v_7004_0 : 3'h0;
  assign v_8333_0 = v_8334_0 | v_8335_0;
  assign v_8334_0 = v_607_0 ? v_7018_0 : 3'h0;
  assign v_8335_0 = v_26_0 ? v_7004_0 : 3'h0;
  assign v_8336_0 = v_601_0 ? v_6997_0 : 3'h0;
  assign v_8337_0 = v_8338_0 | v_8339_0;
  assign v_8338_0 = v_607_0 ? v_7011_0 : 3'h0;
  assign v_8339_0 = v_26_0 ? v_6997_0 : 3'h0;
  assign v_8340_0 = v_601_0 ? v_6990_0 : 3'h0;
  assign v_8341_0 = v_8342_0 | v_8343_0;
  assign v_8342_0 = v_607_0 ? v_7004_0 : 3'h0;
  assign v_8343_0 = v_26_0 ? v_6990_0 : 3'h0;
  assign v_8344_0 = v_601_0 ? v_6983_0 : 3'h0;
  assign v_8345_0 = v_8346_0 | v_8347_0;
  assign v_8346_0 = v_607_0 ? v_6997_0 : 3'h0;
  assign v_8347_0 = v_26_0 ? v_6983_0 : 3'h0;
  assign v_8348_0 = v_601_0 ? v_6976_0 : 3'h0;
  assign v_8349_0 = v_8350_0 | v_8351_0;
  assign v_8350_0 = v_607_0 ? v_6990_0 : 3'h0;
  assign v_8351_0 = v_26_0 ? v_6976_0 : 3'h0;
  assign v_8352_0 = v_601_0 ? v_6969_0 : 3'h0;
  assign v_8353_0 = v_8354_0 | v_8355_0;
  assign v_8354_0 = v_607_0 ? v_6983_0 : 3'h0;
  assign v_8355_0 = v_26_0 ? v_6969_0 : 3'h0;
  assign v_8356_0 = v_601_0 ? v_6962_0 : 3'h0;
  assign v_8357_0 = v_8358_0 | v_8359_0;
  assign v_8358_0 = v_607_0 ? v_6976_0 : 3'h0;
  assign v_8359_0 = v_26_0 ? v_6962_0 : 3'h0;
  assign v_8360_0 = v_601_0 ? v_6955_0 : 3'h0;
  assign v_8361_0 = v_8362_0 | v_8363_0;
  assign v_8362_0 = v_607_0 ? v_6969_0 : 3'h0;
  assign v_8363_0 = v_26_0 ? v_6955_0 : 3'h0;
  assign v_8364_0 = v_601_0 ? v_6948_0 : 3'h0;
  assign v_8365_0 = v_8366_0 | v_8367_0;
  assign v_8366_0 = v_607_0 ? v_6962_0 : 3'h0;
  assign v_8367_0 = v_26_0 ? v_6948_0 : 3'h0;
  assign v_8368_0 = v_601_0 ? v_6941_0 : 3'h0;
  assign v_8369_0 = v_8370_0 | v_8371_0;
  assign v_8370_0 = v_607_0 ? v_6955_0 : 3'h0;
  assign v_8371_0 = v_26_0 ? v_6941_0 : 3'h0;
  assign v_8372_0 = v_601_0 ? v_6934_0 : 3'h0;
  assign v_8373_0 = v_8374_0 | v_8375_0;
  assign v_8374_0 = v_607_0 ? v_6948_0 : 3'h0;
  assign v_8375_0 = v_26_0 ? v_6934_0 : 3'h0;
  assign v_8376_0 = v_601_0 ? v_6927_0 : 3'h0;
  assign v_8377_0 = v_8378_0 | v_8379_0;
  assign v_8378_0 = v_607_0 ? v_6941_0 : 3'h0;
  assign v_8379_0 = v_26_0 ? v_6927_0 : 3'h0;
  assign v_8380_0 = v_601_0 ? v_6920_0 : 3'h0;
  assign v_8381_0 = v_8382_0 | v_8383_0;
  assign v_8382_0 = v_607_0 ? v_6934_0 : 3'h0;
  assign v_8383_0 = v_26_0 ? v_6920_0 : 3'h0;
  assign v_8384_0 = v_601_0 ? v_6913_0 : 3'h0;
  assign v_8385_0 = v_8386_0 | v_8387_0;
  assign v_8386_0 = v_607_0 ? v_6927_0 : 3'h0;
  assign v_8387_0 = v_26_0 ? v_6913_0 : 3'h0;
  assign v_8388_0 = v_601_0 ? v_6906_0 : 3'h0;
  assign v_8389_0 = v_8390_0 | v_8391_0;
  assign v_8390_0 = v_607_0 ? v_6920_0 : 3'h0;
  assign v_8391_0 = v_26_0 ? v_6906_0 : 3'h0;
  assign v_8392_0 = v_601_0 ? v_6899_0 : 3'h0;
  assign v_8393_0 = v_8394_0 | v_8395_0;
  assign v_8394_0 = v_607_0 ? v_6913_0 : 3'h0;
  assign v_8395_0 = v_26_0 ? v_6899_0 : 3'h0;
  assign v_8396_0 = v_601_0 ? v_6892_0 : 3'h0;
  assign v_8397_0 = v_8398_0 | v_8399_0;
  assign v_8398_0 = v_607_0 ? v_6906_0 : 3'h0;
  assign v_8399_0 = v_26_0 ? v_6892_0 : 3'h0;
  assign v_8400_0 = v_601_0 ? v_6885_0 : 3'h0;
  assign v_8401_0 = v_8402_0 | v_8403_0;
  assign v_8402_0 = v_607_0 ? v_6899_0 : 3'h0;
  assign v_8403_0 = v_26_0 ? v_6885_0 : 3'h0;
  assign v_8404_0 = v_601_0 ? v_6878_0 : 3'h0;
  assign v_8405_0 = v_8406_0 | v_8407_0;
  assign v_8406_0 = v_607_0 ? v_6892_0 : 3'h0;
  assign v_8407_0 = v_26_0 ? v_6878_0 : 3'h0;
  assign v_8408_0 = v_601_0 ? v_6871_0 : 3'h0;
  assign v_8409_0 = v_8410_0 | v_8411_0;
  assign v_8410_0 = v_607_0 ? v_6885_0 : 3'h0;
  assign v_8411_0 = v_26_0 ? v_6871_0 : 3'h0;
  assign v_8412_0 = v_601_0 ? v_6864_0 : 3'h0;
  assign v_8413_0 = v_8414_0 | v_8415_0;
  assign v_8414_0 = v_607_0 ? v_6878_0 : 3'h0;
  assign v_8415_0 = v_26_0 ? v_6864_0 : 3'h0;
  assign v_8416_0 = v_601_0 ? v_6857_0 : 3'h0;
  assign v_8417_0 = v_8418_0 | v_8419_0;
  assign v_8418_0 = v_607_0 ? v_6871_0 : 3'h0;
  assign v_8419_0 = v_26_0 ? v_6857_0 : 3'h0;
  assign v_8420_0 = v_601_0 ? v_6850_0 : 3'h0;
  assign v_8421_0 = v_8422_0 | v_8423_0;
  assign v_8422_0 = v_607_0 ? v_6864_0 : 3'h0;
  assign v_8423_0 = v_26_0 ? v_6850_0 : 3'h0;
  assign v_8424_0 = v_601_0 ? v_6843_0 : 3'h0;
  assign v_8425_0 = v_8426_0 | v_8427_0;
  assign v_8426_0 = v_607_0 ? v_6857_0 : 3'h0;
  assign v_8427_0 = v_26_0 ? v_6843_0 : 3'h0;
  assign v_8428_0 = v_601_0 ? v_6836_0 : 3'h0;
  assign v_8429_0 = v_8430_0 | v_8431_0;
  assign v_8430_0 = v_607_0 ? v_6850_0 : 3'h0;
  assign v_8431_0 = v_26_0 ? v_6836_0 : 3'h0;
  assign v_8432_0 = v_601_0 ? v_6829_0 : 3'h0;
  assign v_8433_0 = v_8434_0 | v_8435_0;
  assign v_8434_0 = v_607_0 ? v_6843_0 : 3'h0;
  assign v_8435_0 = v_26_0 ? v_6829_0 : 3'h0;
  assign v_8436_0 = v_601_0 ? v_6822_0 : 3'h0;
  assign v_8437_0 = v_8438_0 | v_8439_0;
  assign v_8438_0 = v_607_0 ? v_6836_0 : 3'h0;
  assign v_8439_0 = v_26_0 ? v_6822_0 : 3'h0;
  assign v_8440_0 = v_601_0 ? v_6815_0 : 3'h0;
  assign v_8441_0 = v_8442_0 | v_8443_0;
  assign v_8442_0 = v_607_0 ? v_6829_0 : 3'h0;
  assign v_8443_0 = v_26_0 ? v_6815_0 : 3'h0;
  assign v_8444_0 = v_601_0 ? v_6808_0 : 3'h0;
  assign v_8445_0 = v_8446_0 | v_8447_0;
  assign v_8446_0 = v_607_0 ? v_6822_0 : 3'h0;
  assign v_8447_0 = v_26_0 ? v_6808_0 : 3'h0;
  assign v_8448_0 = v_601_0 ? v_6801_0 : 3'h0;
  assign v_8449_0 = v_8450_0 | v_8451_0;
  assign v_8450_0 = v_607_0 ? v_6815_0 : 3'h0;
  assign v_8451_0 = v_26_0 ? v_6801_0 : 3'h0;
  assign v_8452_0 = v_601_0 ? v_6794_0 : 3'h0;
  assign v_8453_0 = v_8454_0 | v_8455_0;
  assign v_8454_0 = v_607_0 ? v_6808_0 : 3'h0;
  assign v_8455_0 = v_26_0 ? v_6794_0 : 3'h0;
  assign v_8456_0 = v_601_0 ? v_6787_0 : 3'h0;
  assign v_8457_0 = v_8458_0 | v_8459_0;
  assign v_8458_0 = v_607_0 ? v_6801_0 : 3'h0;
  assign v_8459_0 = v_26_0 ? v_6787_0 : 3'h0;
  assign v_8460_0 = v_601_0 ? v_6780_0 : 3'h0;
  assign v_8461_0 = v_8462_0 | v_8463_0;
  assign v_8462_0 = v_607_0 ? v_6794_0 : 3'h0;
  assign v_8463_0 = v_26_0 ? v_6780_0 : 3'h0;
  assign v_8464_0 = v_601_0 ? v_6773_0 : 3'h0;
  assign v_8465_0 = v_8466_0 | v_8467_0;
  assign v_8466_0 = v_607_0 ? v_6787_0 : 3'h0;
  assign v_8467_0 = v_26_0 ? v_6773_0 : 3'h0;
  assign v_8468_0 = v_601_0 ? v_6766_0 : 3'h0;
  assign v_8469_0 = v_8470_0 | v_8471_0;
  assign v_8470_0 = v_607_0 ? v_6780_0 : 3'h0;
  assign v_8471_0 = v_26_0 ? v_6766_0 : 3'h0;
  assign v_8472_0 = v_601_0 ? v_6759_0 : 3'h0;
  assign v_8473_0 = v_8474_0 | v_8475_0;
  assign v_8474_0 = v_607_0 ? v_6773_0 : 3'h0;
  assign v_8475_0 = v_26_0 ? v_6759_0 : 3'h0;
  assign v_8476_0 = v_601_0 ? v_6752_0 : 3'h0;
  assign v_8477_0 = v_8478_0 | v_8479_0;
  assign v_8478_0 = v_607_0 ? v_6766_0 : 3'h0;
  assign v_8479_0 = v_26_0 ? v_6752_0 : 3'h0;
  assign v_8480_0 = v_601_0 ? v_6745_0 : 3'h0;
  assign v_8481_0 = v_8482_0 | v_8483_0;
  assign v_8482_0 = v_607_0 ? v_6759_0 : 3'h0;
  assign v_8483_0 = v_26_0 ? v_6745_0 : 3'h0;
  assign v_8484_0 = v_601_0 ? v_6738_0 : 3'h0;
  assign v_8485_0 = v_8486_0 | v_8487_0;
  assign v_8486_0 = v_607_0 ? v_6752_0 : 3'h0;
  assign v_8487_0 = v_26_0 ? v_6738_0 : 3'h0;
  assign v_8488_0 = v_601_0 ? v_6731_0 : 3'h0;
  assign v_8489_0 = v_8490_0 | v_8491_0;
  assign v_8490_0 = v_607_0 ? v_6745_0 : 3'h0;
  assign v_8491_0 = v_26_0 ? v_6731_0 : 3'h0;
  assign v_8492_0 = v_601_0 ? v_6724_0 : 3'h0;
  assign v_8493_0 = v_8494_0 | v_8495_0;
  assign v_8494_0 = v_607_0 ? v_6738_0 : 3'h0;
  assign v_8495_0 = v_26_0 ? v_6724_0 : 3'h0;
  assign v_8496_0 = v_601_0 ? v_6717_0 : 3'h0;
  assign v_8497_0 = v_8498_0 | v_8499_0;
  assign v_8498_0 = v_607_0 ? v_6731_0 : 3'h0;
  assign v_8499_0 = v_26_0 ? v_6717_0 : 3'h0;
  assign v_8500_0 = v_601_0 ? v_6710_0 : 3'h0;
  assign v_8501_0 = v_8502_0 | v_8503_0;
  assign v_8502_0 = v_607_0 ? v_6724_0 : 3'h0;
  assign v_8503_0 = v_26_0 ? v_6710_0 : 3'h0;
  assign v_8504_0 = v_601_0 ? v_6703_0 : 3'h0;
  assign v_8505_0 = v_8506_0 | v_8507_0;
  assign v_8506_0 = v_607_0 ? v_6717_0 : 3'h0;
  assign v_8507_0 = v_26_0 ? v_6703_0 : 3'h0;
  assign v_8508_0 = v_601_0 ? v_6696_0 : 3'h0;
  assign v_8509_0 = v_8510_0 | v_8511_0;
  assign v_8510_0 = v_607_0 ? v_6710_0 : 3'h0;
  assign v_8511_0 = v_26_0 ? v_6696_0 : 3'h0;
  assign v_8512_0 = v_601_0 ? v_6689_0 : 3'h0;
  assign v_8513_0 = v_8514_0 | v_8515_0;
  assign v_8514_0 = v_607_0 ? v_6703_0 : 3'h0;
  assign v_8515_0 = v_26_0 ? v_6689_0 : 3'h0;
  assign v_8516_0 = v_601_0 ? v_6682_0 : 3'h0;
  assign v_8517_0 = v_8518_0 | v_8519_0;
  assign v_8518_0 = v_607_0 ? v_6696_0 : 3'h0;
  assign v_8519_0 = v_26_0 ? v_6682_0 : 3'h0;
  assign v_8520_0 = v_601_0 ? v_6675_0 : 3'h0;
  assign v_8521_0 = v_8522_0 | v_8523_0;
  assign v_8522_0 = v_607_0 ? v_6689_0 : 3'h0;
  assign v_8523_0 = v_26_0 ? v_6675_0 : 3'h0;
  assign v_8524_0 = v_601_0 ? v_6668_0 : 3'h0;
  assign v_8525_0 = v_8526_0 | v_8527_0;
  assign v_8526_0 = v_607_0 ? v_6682_0 : 3'h0;
  assign v_8527_0 = v_26_0 ? v_6668_0 : 3'h0;
  assign v_8528_0 = v_601_0 ? v_6661_0 : 3'h0;
  assign v_8529_0 = v_8530_0 | v_8531_0;
  assign v_8530_0 = v_607_0 ? v_6675_0 : 3'h0;
  assign v_8531_0 = v_26_0 ? v_6661_0 : 3'h0;
  assign v_8532_0 = v_601_0 ? v_6654_0 : 3'h0;
  assign v_8533_0 = v_8534_0 | v_8535_0;
  assign v_8534_0 = v_607_0 ? v_6668_0 : 3'h0;
  assign v_8535_0 = v_26_0 ? v_6654_0 : 3'h0;
  assign v_8536_0 = v_601_0 ? v_6647_0 : 3'h0;
  assign v_8537_0 = v_8538_0 | v_8539_0;
  assign v_8538_0 = v_607_0 ? v_6661_0 : 3'h0;
  assign v_8539_0 = v_26_0 ? v_6647_0 : 3'h0;
  assign v_8540_0 = v_601_0 ? v_6640_0 : 3'h0;
  assign v_8541_0 = v_8542_0 | v_8543_0;
  assign v_8542_0 = v_607_0 ? v_6654_0 : 3'h0;
  assign v_8543_0 = v_26_0 ? v_6640_0 : 3'h0;
  assign v_8544_0 = v_601_0 ? v_6633_0 : 3'h0;
  assign v_8545_0 = v_8546_0 | v_8547_0;
  assign v_8546_0 = v_607_0 ? v_6647_0 : 3'h0;
  assign v_8547_0 = v_26_0 ? v_6633_0 : 3'h0;
  assign v_8548_0 = v_601_0 ? v_6626_0 : 3'h0;
  assign v_8549_0 = v_8550_0 | v_8551_0;
  assign v_8550_0 = v_607_0 ? v_6640_0 : 3'h0;
  assign v_8551_0 = v_26_0 ? v_6626_0 : 3'h0;
  assign v_8552_0 = v_601_0 ? v_6619_0 : 3'h0;
  assign v_8553_0 = v_8554_0 | v_8555_0;
  assign v_8554_0 = v_607_0 ? v_6633_0 : 3'h0;
  assign v_8555_0 = v_26_0 ? v_6619_0 : 3'h0;
  assign v_8556_0 = v_601_0 ? v_6612_0 : 3'h0;
  assign v_8557_0 = v_8558_0 | v_8559_0;
  assign v_8558_0 = v_607_0 ? v_6626_0 : 3'h0;
  assign v_8559_0 = v_26_0 ? v_6612_0 : 3'h0;
  assign v_8560_0 = v_601_0 ? v_6605_0 : 3'h0;
  assign v_8561_0 = v_8562_0 | v_8563_0;
  assign v_8562_0 = v_607_0 ? v_6619_0 : 3'h0;
  assign v_8563_0 = v_26_0 ? v_6605_0 : 3'h0;
  assign v_8564_0 = v_601_0 ? v_6598_0 : 3'h0;
  assign v_8565_0 = v_8566_0 | v_8567_0;
  assign v_8566_0 = v_607_0 ? v_6612_0 : 3'h0;
  assign v_8567_0 = v_26_0 ? v_6598_0 : 3'h0;
  assign v_8568_0 = v_601_0 ? v_6591_0 : 3'h0;
  assign v_8569_0 = v_8570_0 | v_8571_0;
  assign v_8570_0 = v_607_0 ? v_6605_0 : 3'h0;
  assign v_8571_0 = v_26_0 ? v_6591_0 : 3'h0;
  assign v_8572_0 = v_601_0 ? v_6584_0 : 3'h0;
  assign v_8573_0 = v_8574_0 | v_8575_0;
  assign v_8574_0 = v_607_0 ? v_6598_0 : 3'h0;
  assign v_8575_0 = v_26_0 ? v_6584_0 : 3'h0;
  assign v_8576_0 = v_601_0 ? v_6577_0 : 3'h0;
  assign v_8577_0 = v_8578_0 | v_8579_0;
  assign v_8578_0 = v_607_0 ? v_6591_0 : 3'h0;
  assign v_8579_0 = v_26_0 ? v_6577_0 : 3'h0;
  assign v_8580_0 = v_601_0 ? v_6570_0 : 3'h0;
  assign v_8581_0 = v_8582_0 | v_8583_0;
  assign v_8582_0 = v_607_0 ? v_6584_0 : 3'h0;
  assign v_8583_0 = v_26_0 ? v_6570_0 : 3'h0;
  assign v_8584_0 = v_601_0 ? v_6563_0 : 3'h0;
  assign v_8585_0 = v_8586_0 | v_8587_0;
  assign v_8586_0 = v_607_0 ? v_6577_0 : 3'h0;
  assign v_8587_0 = v_26_0 ? v_6563_0 : 3'h0;
  assign v_8588_0 = v_601_0 ? v_6556_0 : 3'h0;
  assign v_8589_0 = v_8590_0 | v_8591_0;
  assign v_8590_0 = v_607_0 ? v_6570_0 : 3'h0;
  assign v_8591_0 = v_26_0 ? v_6556_0 : 3'h0;
  assign v_8592_0 = v_601_0 ? v_6549_0 : 3'h0;
  assign v_8593_0 = v_8594_0 | v_8595_0;
  assign v_8594_0 = v_607_0 ? v_6563_0 : 3'h0;
  assign v_8595_0 = v_26_0 ? v_6549_0 : 3'h0;
  assign v_8596_0 = v_601_0 ? v_6542_0 : 3'h0;
  assign v_8597_0 = v_8598_0 | v_8599_0;
  assign v_8598_0 = v_607_0 ? v_6556_0 : 3'h0;
  assign v_8599_0 = v_26_0 ? v_6542_0 : 3'h0;
  assign v_8600_0 = v_601_0 ? v_6535_0 : 3'h0;
  assign v_8601_0 = v_8602_0 | v_8603_0;
  assign v_8602_0 = v_607_0 ? v_6549_0 : 3'h0;
  assign v_8603_0 = v_26_0 ? v_6535_0 : 3'h0;
  assign v_8604_0 = v_601_0 ? v_6528_0 : 3'h0;
  assign v_8605_0 = v_8606_0 | v_8607_0;
  assign v_8606_0 = v_607_0 ? v_6542_0 : 3'h0;
  assign v_8607_0 = v_26_0 ? v_6528_0 : 3'h0;
  assign v_8608_0 = v_601_0 ? v_6521_0 : 3'h0;
  assign v_8609_0 = v_8610_0 | v_8611_0;
  assign v_8610_0 = v_607_0 ? v_6535_0 : 3'h0;
  assign v_8611_0 = v_26_0 ? v_6521_0 : 3'h0;
  assign v_8612_0 = v_601_0 ? v_6514_0 : 3'h0;
  assign v_8613_0 = v_8614_0 | v_8615_0;
  assign v_8614_0 = v_607_0 ? v_6528_0 : 3'h0;
  assign v_8615_0 = v_26_0 ? v_6514_0 : 3'h0;
  assign v_8616_0 = v_601_0 ? v_6507_0 : 3'h0;
  assign v_8617_0 = v_8618_0 | v_8619_0;
  assign v_8618_0 = v_607_0 ? v_6521_0 : 3'h0;
  assign v_8619_0 = v_26_0 ? v_6507_0 : 3'h0;
  assign v_8620_0 = v_601_0 ? v_6500_0 : 3'h0;
  assign v_8621_0 = v_8622_0 | v_8623_0;
  assign v_8622_0 = v_607_0 ? v_6514_0 : 3'h0;
  assign v_8623_0 = v_26_0 ? v_6500_0 : 3'h0;
  assign v_8624_0 = v_601_0 ? v_6493_0 : 3'h0;
  assign v_8625_0 = v_8626_0 | v_8627_0;
  assign v_8626_0 = v_607_0 ? v_6507_0 : 3'h0;
  assign v_8627_0 = v_26_0 ? v_6493_0 : 3'h0;
  assign v_8628_0 = v_601_0 ? v_6486_0 : 3'h0;
  assign v_8629_0 = v_8630_0 | v_8631_0;
  assign v_8630_0 = v_607_0 ? v_6500_0 : 3'h0;
  assign v_8631_0 = v_26_0 ? v_6486_0 : 3'h0;
  assign v_8632_0 = v_601_0 ? v_6479_0 : 3'h0;
  assign v_8633_0 = v_8634_0 | v_8635_0;
  assign v_8634_0 = v_607_0 ? v_6493_0 : 3'h0;
  assign v_8635_0 = v_26_0 ? v_6479_0 : 3'h0;
  assign v_8636_0 = v_601_0 ? v_6472_0 : 3'h0;
  assign v_8637_0 = v_8638_0 | v_8639_0;
  assign v_8638_0 = v_607_0 ? v_6486_0 : 3'h0;
  assign v_8639_0 = v_26_0 ? v_6472_0 : 3'h0;
  assign v_8640_0 = v_601_0 ? v_6465_0 : 3'h0;
  assign v_8641_0 = v_8642_0 | v_8643_0;
  assign v_8642_0 = v_607_0 ? v_6479_0 : 3'h0;
  assign v_8643_0 = v_26_0 ? v_6465_0 : 3'h0;
  assign v_8644_0 = v_601_0 ? v_6458_0 : 3'h0;
  assign v_8645_0 = v_8646_0 | v_8647_0;
  assign v_8646_0 = v_607_0 ? v_6472_0 : 3'h0;
  assign v_8647_0 = v_26_0 ? v_6458_0 : 3'h0;
  assign v_8648_0 = v_601_0 ? v_6451_0 : 3'h0;
  assign v_8649_0 = v_8650_0 | v_8651_0;
  assign v_8650_0 = v_607_0 ? v_6465_0 : 3'h0;
  assign v_8651_0 = v_26_0 ? v_6451_0 : 3'h0;
  assign v_8652_0 = v_601_0 ? v_6444_0 : 3'h0;
  assign v_8653_0 = v_8654_0 | v_8655_0;
  assign v_8654_0 = v_607_0 ? v_6458_0 : 3'h0;
  assign v_8655_0 = v_26_0 ? v_6444_0 : 3'h0;
  assign v_8656_0 = v_601_0 ? v_6437_0 : 3'h0;
  assign v_8657_0 = v_8658_0 | v_8659_0;
  assign v_8658_0 = v_607_0 ? v_6451_0 : 3'h0;
  assign v_8659_0 = v_26_0 ? v_6437_0 : 3'h0;
  assign v_8660_0 = v_601_0 ? v_6430_0 : 3'h0;
  assign v_8661_0 = v_8662_0 | v_8663_0;
  assign v_8662_0 = v_607_0 ? v_6444_0 : 3'h0;
  assign v_8663_0 = v_26_0 ? v_6430_0 : 3'h0;
  assign v_8664_0 = v_601_0 ? v_6423_0 : 3'h0;
  assign v_8665_0 = v_8666_0 | v_8667_0;
  assign v_8666_0 = v_607_0 ? v_6437_0 : 3'h0;
  assign v_8667_0 = v_26_0 ? v_6423_0 : 3'h0;
  assign v_8668_0 = v_601_0 ? v_6416_0 : 3'h0;
  assign v_8669_0 = v_8670_0 | v_8671_0;
  assign v_8670_0 = v_607_0 ? v_6430_0 : 3'h0;
  assign v_8671_0 = v_26_0 ? v_6416_0 : 3'h0;
  assign v_8672_0 = v_601_0 ? v_6409_0 : 3'h0;
  assign v_8673_0 = v_8674_0 | v_8675_0;
  assign v_8674_0 = v_607_0 ? v_6423_0 : 3'h0;
  assign v_8675_0 = v_26_0 ? v_6409_0 : 3'h0;
  assign v_8676_0 = v_601_0 ? v_6402_0 : 3'h0;
  assign v_8677_0 = v_8678_0 | v_8679_0;
  assign v_8678_0 = v_607_0 ? v_6416_0 : 3'h0;
  assign v_8679_0 = v_26_0 ? v_6402_0 : 3'h0;
  assign v_8680_0 = v_601_0 ? v_6395_0 : 3'h0;
  assign v_8681_0 = v_8682_0 | v_8683_0;
  assign v_8682_0 = v_607_0 ? v_6409_0 : 3'h0;
  assign v_8683_0 = v_26_0 ? v_6395_0 : 3'h0;
  assign v_8684_0 = v_601_0 ? v_6388_0 : 3'h0;
  assign v_8685_0 = v_8686_0 | v_8687_0;
  assign v_8686_0 = v_607_0 ? v_6402_0 : 3'h0;
  assign v_8687_0 = v_26_0 ? v_6388_0 : 3'h0;
  assign v_8688_0 = v_601_0 ? v_6381_0 : 3'h0;
  assign v_8689_0 = v_8690_0 | v_8691_0;
  assign v_8690_0 = v_607_0 ? v_6395_0 : 3'h0;
  assign v_8691_0 = v_26_0 ? v_6381_0 : 3'h0;
  assign v_8692_0 = v_601_0 ? v_6374_0 : 3'h0;
  assign v_8693_0 = v_8694_0 | v_8695_0;
  assign v_8694_0 = v_607_0 ? v_6388_0 : 3'h0;
  assign v_8695_0 = v_26_0 ? v_6374_0 : 3'h0;
  assign v_8696_0 = v_601_0 ? v_6367_0 : 3'h0;
  assign v_8697_0 = v_8698_0 | v_8699_0;
  assign v_8698_0 = v_607_0 ? v_6381_0 : 3'h0;
  assign v_8699_0 = v_26_0 ? v_6367_0 : 3'h0;
  assign v_8700_0 = v_601_0 ? v_6360_0 : 3'h0;
  assign v_8701_0 = v_8702_0 | v_8703_0;
  assign v_8702_0 = v_607_0 ? v_6374_0 : 3'h0;
  assign v_8703_0 = v_26_0 ? v_6360_0 : 3'h0;
  assign v_8704_0 = v_601_0 ? v_6353_0 : 3'h0;
  assign v_8705_0 = v_8706_0 | v_8707_0;
  assign v_8706_0 = v_607_0 ? v_6367_0 : 3'h0;
  assign v_8707_0 = v_26_0 ? v_6353_0 : 3'h0;
  assign v_8708_0 = v_601_0 ? v_6346_0 : 3'h0;
  assign v_8709_0 = v_8710_0 | v_8711_0;
  assign v_8710_0 = v_607_0 ? v_6360_0 : 3'h0;
  assign v_8711_0 = v_26_0 ? v_6346_0 : 3'h0;
  assign v_8712_0 = v_601_0 ? v_6339_0 : 3'h0;
  assign v_8713_0 = v_8714_0 | v_8715_0;
  assign v_8714_0 = v_607_0 ? v_6353_0 : 3'h0;
  assign v_8715_0 = v_26_0 ? v_6339_0 : 3'h0;
  assign v_8716_0 = v_601_0 ? v_6332_0 : 3'h0;
  assign v_8717_0 = v_8718_0 | v_8719_0;
  assign v_8718_0 = v_607_0 ? v_6346_0 : 3'h0;
  assign v_8719_0 = v_26_0 ? v_6332_0 : 3'h0;
  assign v_8720_0 = v_601_0 ? v_6325_0 : 3'h0;
  assign v_8721_0 = v_8722_0 | v_8723_0;
  assign v_8722_0 = v_607_0 ? v_6339_0 : 3'h0;
  assign v_8723_0 = v_26_0 ? v_6325_0 : 3'h0;
  assign v_8724_0 = v_601_0 ? v_6318_0 : 3'h0;
  assign v_8725_0 = v_8726_0 | v_8727_0;
  assign v_8726_0 = v_607_0 ? v_6332_0 : 3'h0;
  assign v_8727_0 = v_26_0 ? v_6318_0 : 3'h0;
  assign v_8728_0 = v_601_0 ? v_6311_0 : 3'h0;
  assign v_8729_0 = v_8730_0 | v_8731_0;
  assign v_8730_0 = v_607_0 ? v_6325_0 : 3'h0;
  assign v_8731_0 = v_26_0 ? v_6311_0 : 3'h0;
  assign v_8732_0 = v_601_0 ? v_6304_0 : 3'h0;
  assign v_8733_0 = v_8734_0 | v_8735_0;
  assign v_8734_0 = v_607_0 ? v_6318_0 : 3'h0;
  assign v_8735_0 = v_26_0 ? v_6304_0 : 3'h0;
  assign v_8736_0 = v_601_0 ? v_6297_0 : 3'h0;
  assign v_8737_0 = v_8738_0 | v_8739_0;
  assign v_8738_0 = v_607_0 ? v_6311_0 : 3'h0;
  assign v_8739_0 = v_26_0 ? v_6297_0 : 3'h0;
  assign v_8740_0 = v_601_0 ? v_6290_0 : 3'h0;
  assign v_8741_0 = v_8742_0 | v_8743_0;
  assign v_8742_0 = v_607_0 ? v_6304_0 : 3'h0;
  assign v_8743_0 = v_26_0 ? v_6290_0 : 3'h0;
  assign v_8744_0 = v_601_0 ? v_6283_0 : 3'h0;
  assign v_8745_0 = v_8746_0 | v_8747_0;
  assign v_8746_0 = v_607_0 ? v_6297_0 : 3'h0;
  assign v_8747_0 = v_26_0 ? v_6283_0 : 3'h0;
  assign v_8748_0 = v_601_0 ? v_6276_0 : 3'h0;
  assign v_8749_0 = v_8750_0 | v_8751_0;
  assign v_8750_0 = v_607_0 ? v_6290_0 : 3'h0;
  assign v_8751_0 = v_26_0 ? v_6276_0 : 3'h0;
  assign v_8752_0 = v_601_0 ? v_6269_0 : 3'h0;
  assign v_8753_0 = v_8754_0 | v_8755_0;
  assign v_8754_0 = v_607_0 ? v_6283_0 : 3'h0;
  assign v_8755_0 = v_26_0 ? v_6269_0 : 3'h0;
  assign v_8756_0 = v_601_0 ? v_6262_0 : 3'h0;
  assign v_8757_0 = v_8758_0 | v_8759_0;
  assign v_8758_0 = v_607_0 ? v_6276_0 : 3'h0;
  assign v_8759_0 = v_26_0 ? v_6262_0 : 3'h0;
  assign v_8760_0 = v_601_0 ? v_6255_0 : 3'h0;
  assign v_8761_0 = v_8762_0 | v_8763_0;
  assign v_8762_0 = v_607_0 ? v_6269_0 : 3'h0;
  assign v_8763_0 = v_26_0 ? v_6255_0 : 3'h0;
  assign v_8764_0 = v_601_0 ? v_6248_0 : 3'h0;
  assign v_8765_0 = v_8766_0 | v_8767_0;
  assign v_8766_0 = v_607_0 ? v_6262_0 : 3'h0;
  assign v_8767_0 = v_26_0 ? v_6248_0 : 3'h0;
  assign v_8768_0 = v_601_0 ? v_6241_0 : 3'h0;
  assign v_8769_0 = v_8770_0 | v_8771_0;
  assign v_8770_0 = v_607_0 ? v_6255_0 : 3'h0;
  assign v_8771_0 = v_26_0 ? v_6241_0 : 3'h0;
  assign v_8772_0 = v_601_0 ? v_6234_0 : 3'h0;
  assign v_8773_0 = v_8774_0 | v_8775_0;
  assign v_8774_0 = v_607_0 ? v_6248_0 : 3'h0;
  assign v_8775_0 = v_26_0 ? v_6234_0 : 3'h0;
  assign v_8776_0 = v_601_0 ? v_6227_0 : 3'h0;
  assign v_8777_0 = v_8778_0 | v_8779_0;
  assign v_8778_0 = v_607_0 ? v_6241_0 : 3'h0;
  assign v_8779_0 = v_26_0 ? v_6227_0 : 3'h0;
  assign v_8780_0 = v_601_0 ? v_6220_0 : 3'h0;
  assign v_8781_0 = v_8782_0 | v_8783_0;
  assign v_8782_0 = v_607_0 ? v_6234_0 : 3'h0;
  assign v_8783_0 = v_26_0 ? v_6220_0 : 3'h0;
  assign v_8784_0 = v_601_0 ? v_6213_0 : 3'h0;
  assign v_8785_0 = v_8786_0 | v_8787_0;
  assign v_8786_0 = v_607_0 ? v_6227_0 : 3'h0;
  assign v_8787_0 = v_26_0 ? v_6213_0 : 3'h0;
  assign v_8788_0 = v_601_0 ? v_6206_0 : 3'h0;
  assign v_8789_0 = v_8790_0 | v_8791_0;
  assign v_8790_0 = v_607_0 ? v_6220_0 : 3'h0;
  assign v_8791_0 = v_26_0 ? v_6206_0 : 3'h0;
  assign v_8792_0 = v_601_0 ? v_6199_0 : 3'h0;
  assign v_8793_0 = v_8794_0 | v_8795_0;
  assign v_8794_0 = v_607_0 ? v_6213_0 : 3'h0;
  assign v_8795_0 = v_26_0 ? v_6199_0 : 3'h0;
  assign v_8796_0 = v_601_0 ? v_6192_0 : 3'h0;
  assign v_8797_0 = v_8798_0 | v_8799_0;
  assign v_8798_0 = v_607_0 ? v_6206_0 : 3'h0;
  assign v_8799_0 = v_26_0 ? v_6192_0 : 3'h0;
  assign v_8800_0 = v_601_0 ? v_6185_0 : 3'h0;
  assign v_8801_0 = v_8802_0 | v_8803_0;
  assign v_8802_0 = v_607_0 ? v_6199_0 : 3'h0;
  assign v_8803_0 = v_26_0 ? v_6185_0 : 3'h0;
  assign v_8804_0 = v_601_0 ? v_6178_0 : 3'h0;
  assign v_8805_0 = v_8806_0 | v_8807_0;
  assign v_8806_0 = v_607_0 ? v_6192_0 : 3'h0;
  assign v_8807_0 = v_26_0 ? v_6178_0 : 3'h0;
  assign v_8808_0 = v_601_0 ? v_6171_0 : 3'h0;
  assign v_8809_0 = v_8810_0 | v_8811_0;
  assign v_8810_0 = v_607_0 ? v_6185_0 : 3'h0;
  assign v_8811_0 = v_26_0 ? v_6171_0 : 3'h0;
  assign v_8812_0 = v_601_0 ? v_6164_0 : 3'h0;
  assign v_8813_0 = v_8814_0 | v_8815_0;
  assign v_8814_0 = v_607_0 ? v_6178_0 : 3'h0;
  assign v_8815_0 = v_26_0 ? v_6164_0 : 3'h0;
  assign v_8816_0 = v_601_0 ? v_6157_0 : 3'h0;
  assign v_8817_0 = v_8818_0 | v_8819_0;
  assign v_8818_0 = v_607_0 ? v_6171_0 : 3'h0;
  assign v_8819_0 = v_26_0 ? v_6157_0 : 3'h0;
  assign v_8820_0 = v_601_0 ? v_6150_0 : 3'h0;
  assign v_8821_0 = v_8822_0 | v_8823_0;
  assign v_8822_0 = v_607_0 ? v_6164_0 : 3'h0;
  assign v_8823_0 = v_26_0 ? v_6150_0 : 3'h0;
  assign v_8824_0 = v_601_0 ? v_6143_0 : 3'h0;
  assign v_8825_0 = v_8826_0 | v_8827_0;
  assign v_8826_0 = v_607_0 ? v_6157_0 : 3'h0;
  assign v_8827_0 = v_26_0 ? v_6143_0 : 3'h0;
  assign v_8828_0 = v_601_0 ? v_6136_0 : 3'h0;
  assign v_8829_0 = v_8830_0 | v_8831_0;
  assign v_8830_0 = v_607_0 ? v_6150_0 : 3'h0;
  assign v_8831_0 = v_26_0 ? v_6136_0 : 3'h0;
  assign v_8832_0 = v_601_0 ? v_6129_0 : 3'h0;
  assign v_8833_0 = v_8834_0 | v_8835_0;
  assign v_8834_0 = v_607_0 ? v_6143_0 : 3'h0;
  assign v_8835_0 = v_26_0 ? v_6129_0 : 3'h0;
  assign v_8836_0 = v_601_0 ? v_6122_0 : 3'h0;
  assign v_8837_0 = v_8838_0 | v_8839_0;
  assign v_8838_0 = v_607_0 ? v_6136_0 : 3'h0;
  assign v_8839_0 = v_26_0 ? v_6122_0 : 3'h0;
  assign v_8840_0 = v_601_0 ? v_6115_0 : 3'h0;
  assign v_8841_0 = v_8842_0 | v_8843_0;
  assign v_8842_0 = v_607_0 ? v_6129_0 : 3'h0;
  assign v_8843_0 = v_26_0 ? v_6115_0 : 3'h0;
  assign v_8844_0 = v_601_0 ? v_6108_0 : 3'h0;
  assign v_8845_0 = v_8846_0 | v_8847_0;
  assign v_8846_0 = v_607_0 ? v_6122_0 : 3'h0;
  assign v_8847_0 = v_26_0 ? v_6108_0 : 3'h0;
  assign v_8848_0 = v_601_0 ? v_6101_0 : 3'h0;
  assign v_8849_0 = v_8850_0 | v_8851_0;
  assign v_8850_0 = v_607_0 ? v_6115_0 : 3'h0;
  assign v_8851_0 = v_26_0 ? v_6101_0 : 3'h0;
  assign v_8852_0 = v_601_0 ? v_6094_0 : 3'h0;
  assign v_8853_0 = v_8854_0 | v_8855_0;
  assign v_8854_0 = v_607_0 ? v_6108_0 : 3'h0;
  assign v_8855_0 = v_26_0 ? v_6094_0 : 3'h0;
  assign v_8856_0 = v_601_0 ? v_6087_0 : 3'h0;
  assign v_8857_0 = v_8858_0 | v_8859_0;
  assign v_8858_0 = v_607_0 ? v_6101_0 : 3'h0;
  assign v_8859_0 = v_26_0 ? v_6087_0 : 3'h0;
  assign v_8860_0 = v_601_0 ? v_6080_0 : 3'h0;
  assign v_8861_0 = v_8862_0 | v_8863_0;
  assign v_8862_0 = v_607_0 ? v_6094_0 : 3'h0;
  assign v_8863_0 = v_26_0 ? v_6080_0 : 3'h0;
  assign v_8864_0 = v_601_0 ? v_6073_0 : 3'h0;
  assign v_8865_0 = v_8866_0 | v_8867_0;
  assign v_8866_0 = v_607_0 ? v_6087_0 : 3'h0;
  assign v_8867_0 = v_26_0 ? v_6073_0 : 3'h0;
  assign v_8868_0 = v_601_0 ? v_6066_0 : 3'h0;
  assign v_8869_0 = v_8870_0 | v_8871_0;
  assign v_8870_0 = v_607_0 ? v_6080_0 : 3'h0;
  assign v_8871_0 = v_26_0 ? v_6066_0 : 3'h0;
  assign v_8872_0 = v_601_0 ? v_6059_0 : 3'h0;
  assign v_8873_0 = v_8874_0 | v_8875_0;
  assign v_8874_0 = v_607_0 ? v_6073_0 : 3'h0;
  assign v_8875_0 = v_26_0 ? v_6059_0 : 3'h0;
  assign v_8876_0 = v_601_0 ? v_6052_0 : 3'h0;
  assign v_8877_0 = v_8878_0 | v_8879_0;
  assign v_8878_0 = v_607_0 ? v_6066_0 : 3'h0;
  assign v_8879_0 = v_26_0 ? v_6052_0 : 3'h0;
  assign v_8880_0 = v_601_0 ? v_6045_0 : 3'h0;
  assign v_8881_0 = v_8882_0 | v_8883_0;
  assign v_8882_0 = v_607_0 ? v_6059_0 : 3'h0;
  assign v_8883_0 = v_26_0 ? v_6045_0 : 3'h0;
  assign v_8884_0 = v_601_0 ? v_6038_0 : 3'h0;
  assign v_8885_0 = v_8886_0 | v_8887_0;
  assign v_8886_0 = v_607_0 ? v_6052_0 : 3'h0;
  assign v_8887_0 = v_26_0 ? v_6038_0 : 3'h0;
  assign v_8888_0 = v_601_0 ? v_6031_0 : 3'h0;
  assign v_8889_0 = v_8890_0 | v_8891_0;
  assign v_8890_0 = v_607_0 ? v_6045_0 : 3'h0;
  assign v_8891_0 = v_26_0 ? v_6031_0 : 3'h0;
  assign v_8892_0 = v_601_0 ? v_6024_0 : 3'h0;
  assign v_8893_0 = v_8894_0 | v_8895_0;
  assign v_8894_0 = v_607_0 ? v_6038_0 : 3'h0;
  assign v_8895_0 = v_26_0 ? v_6024_0 : 3'h0;
  assign v_8896_0 = v_601_0 ? v_6017_0 : 3'h0;
  assign v_8897_0 = v_8898_0 | v_8899_0;
  assign v_8898_0 = v_607_0 ? v_6031_0 : 3'h0;
  assign v_8899_0 = v_26_0 ? v_6017_0 : 3'h0;
  assign v_8900_0 = v_601_0 ? v_6010_0 : 3'h0;
  assign v_8901_0 = v_8902_0 | v_8903_0;
  assign v_8902_0 = v_607_0 ? v_6024_0 : 3'h0;
  assign v_8903_0 = v_26_0 ? v_6010_0 : 3'h0;
  assign v_8904_0 = v_601_0 ? v_6003_0 : 3'h0;
  assign v_8905_0 = v_8906_0 | v_8907_0;
  assign v_8906_0 = v_607_0 ? v_6017_0 : 3'h0;
  assign v_8907_0 = v_26_0 ? v_6003_0 : 3'h0;
  assign v_8908_0 = v_601_0 ? v_5996_0 : 3'h0;
  assign v_8909_0 = v_8910_0 | v_8911_0;
  assign v_8910_0 = v_607_0 ? v_6010_0 : 3'h0;
  assign v_8911_0 = v_26_0 ? v_5996_0 : 3'h0;
  assign v_8912_0 = v_601_0 ? v_5989_0 : 3'h0;
  assign v_8913_0 = v_8914_0 | v_8915_0;
  assign v_8914_0 = v_607_0 ? v_6003_0 : 3'h0;
  assign v_8915_0 = v_26_0 ? v_5989_0 : 3'h0;
  assign v_8916_0 = v_601_0 ? v_5982_0 : 3'h0;
  assign v_8917_0 = v_8918_0 | v_8919_0;
  assign v_8918_0 = v_607_0 ? v_5996_0 : 3'h0;
  assign v_8919_0 = v_26_0 ? v_5982_0 : 3'h0;
  assign v_8920_0 = v_601_0 ? v_5975_0 : 3'h0;
  assign v_8921_0 = v_8922_0 | v_8923_0;
  assign v_8922_0 = v_607_0 ? v_5989_0 : 3'h0;
  assign v_8923_0 = v_26_0 ? v_5975_0 : 3'h0;
  assign v_8924_0 = v_601_0 ? v_5968_0 : 3'h0;
  assign v_8925_0 = v_8926_0 | v_8927_0;
  assign v_8926_0 = v_607_0 ? v_5982_0 : 3'h0;
  assign v_8927_0 = v_26_0 ? v_5968_0 : 3'h0;
  assign v_8928_0 = v_601_0 ? v_5961_0 : 3'h0;
  assign v_8929_0 = v_8930_0 | v_8931_0;
  assign v_8930_0 = v_607_0 ? v_5975_0 : 3'h0;
  assign v_8931_0 = v_26_0 ? v_5961_0 : 3'h0;
  assign v_8932_0 = v_601_0 ? v_5954_0 : 3'h0;
  assign v_8933_0 = v_8934_0 | v_8935_0;
  assign v_8934_0 = v_607_0 ? v_5968_0 : 3'h0;
  assign v_8935_0 = v_26_0 ? v_5954_0 : 3'h0;
  assign v_8936_0 = v_601_0 ? v_5947_0 : 3'h0;
  assign v_8937_0 = v_8938_0 | v_8939_0;
  assign v_8938_0 = v_607_0 ? v_5961_0 : 3'h0;
  assign v_8939_0 = v_26_0 ? v_5947_0 : 3'h0;
  assign v_8940_0 = v_601_0 ? v_5940_0 : 3'h0;
  assign v_8941_0 = v_8942_0 | v_8943_0;
  assign v_8942_0 = v_607_0 ? v_5954_0 : 3'h0;
  assign v_8943_0 = v_26_0 ? v_5940_0 : 3'h0;
  assign v_8944_0 = v_601_0 ? v_5933_0 : 3'h0;
  assign v_8945_0 = v_8946_0 | v_8947_0;
  assign v_8946_0 = v_607_0 ? v_5947_0 : 3'h0;
  assign v_8947_0 = v_26_0 ? v_5933_0 : 3'h0;
  assign v_8948_0 = v_601_0 ? v_5926_0 : 3'h0;
  assign v_8949_0 = v_8950_0 | v_8951_0;
  assign v_8950_0 = v_607_0 ? v_5940_0 : 3'h0;
  assign v_8951_0 = v_26_0 ? v_5926_0 : 3'h0;
  assign v_8952_0 = v_601_0 ? v_5919_0 : 3'h0;
  assign v_8953_0 = v_8954_0 | v_8955_0;
  assign v_8954_0 = v_607_0 ? v_5933_0 : 3'h0;
  assign v_8955_0 = v_26_0 ? v_5919_0 : 3'h0;
  assign v_8956_0 = v_601_0 ? v_5912_0 : 3'h0;
  assign v_8957_0 = v_8958_0 | v_8959_0;
  assign v_8958_0 = v_607_0 ? v_5926_0 : 3'h0;
  assign v_8959_0 = v_26_0 ? v_5912_0 : 3'h0;
  assign v_8960_0 = v_601_0 ? v_5905_0 : 3'h0;
  assign v_8961_0 = v_8962_0 | v_8963_0;
  assign v_8962_0 = v_607_0 ? v_5919_0 : 3'h0;
  assign v_8963_0 = v_26_0 ? v_5905_0 : 3'h0;
  assign v_8964_0 = v_601_0 ? v_5898_0 : 3'h0;
  assign v_8965_0 = v_8966_0 | v_8967_0;
  assign v_8966_0 = v_607_0 ? v_5912_0 : 3'h0;
  assign v_8967_0 = v_26_0 ? v_5898_0 : 3'h0;
  assign v_8968_0 = v_601_0 ? v_5891_0 : 3'h0;
  assign v_8969_0 = v_8970_0 | v_8971_0;
  assign v_8970_0 = v_607_0 ? v_5905_0 : 3'h0;
  assign v_8971_0 = v_26_0 ? v_5891_0 : 3'h0;
  assign v_8972_0 = v_601_0 ? v_5884_0 : 3'h0;
  assign v_8973_0 = v_8974_0 | v_8975_0;
  assign v_8974_0 = v_607_0 ? v_5898_0 : 3'h0;
  assign v_8975_0 = v_26_0 ? v_5884_0 : 3'h0;
  assign v_8976_0 = v_601_0 ? v_5877_0 : 3'h0;
  assign v_8977_0 = v_8978_0 | v_8979_0;
  assign v_8978_0 = v_607_0 ? v_5891_0 : 3'h0;
  assign v_8979_0 = v_26_0 ? v_5877_0 : 3'h0;
  assign v_8980_0 = v_601_0 ? v_5870_0 : 3'h0;
  assign v_8981_0 = v_8982_0 | v_8983_0;
  assign v_8982_0 = v_607_0 ? v_5884_0 : 3'h0;
  assign v_8983_0 = v_26_0 ? v_5870_0 : 3'h0;
  assign v_8984_0 = v_601_0 ? v_5863_0 : 3'h0;
  assign v_8985_0 = v_8986_0 | v_8987_0;
  assign v_8986_0 = v_607_0 ? v_5877_0 : 3'h0;
  assign v_8987_0 = v_26_0 ? v_5863_0 : 3'h0;
  assign v_8988_0 = v_601_0 ? v_5856_0 : 3'h0;
  assign v_8989_0 = v_8990_0 | v_8991_0;
  assign v_8990_0 = v_607_0 ? v_5870_0 : 3'h0;
  assign v_8991_0 = v_26_0 ? v_5856_0 : 3'h0;
  assign v_8992_0 = v_601_0 ? v_5849_0 : 3'h0;
  assign v_8993_0 = v_8994_0 | v_8995_0;
  assign v_8994_0 = v_607_0 ? v_5863_0 : 3'h0;
  assign v_8995_0 = v_26_0 ? v_5849_0 : 3'h0;
  assign v_8996_0 = v_601_0 ? v_5842_0 : 3'h0;
  assign v_8997_0 = v_8998_0 | v_8999_0;
  assign v_8998_0 = v_607_0 ? v_5856_0 : 3'h0;
  assign v_8999_0 = v_26_0 ? v_5842_0 : 3'h0;
  assign v_9000_0 = v_601_0 ? v_5835_0 : 3'h0;
  assign v_9001_0 = v_9002_0 | v_9003_0;
  assign v_9002_0 = v_607_0 ? v_5849_0 : 3'h0;
  assign v_9003_0 = v_26_0 ? v_5835_0 : 3'h0;
  assign v_9004_0 = v_601_0 ? v_5828_0 : 3'h0;
  assign v_9005_0 = v_9006_0 | v_9007_0;
  assign v_9006_0 = v_607_0 ? v_5842_0 : 3'h0;
  assign v_9007_0 = v_26_0 ? v_5828_0 : 3'h0;
  assign v_9008_0 = v_601_0 ? v_5821_0 : 3'h0;
  assign v_9009_0 = v_9010_0 | v_9011_0;
  assign v_9010_0 = v_607_0 ? v_5835_0 : 3'h0;
  assign v_9011_0 = v_26_0 ? v_5821_0 : 3'h0;
  assign v_9012_0 = v_601_0 ? v_5814_0 : 3'h0;
  assign v_9013_0 = v_9014_0 | v_9015_0;
  assign v_9014_0 = v_607_0 ? v_5828_0 : 3'h0;
  assign v_9015_0 = v_26_0 ? v_5814_0 : 3'h0;
  assign v_9016_0 = v_601_0 ? v_5807_0 : 3'h0;
  assign v_9017_0 = v_9018_0 | v_9019_0;
  assign v_9018_0 = v_607_0 ? v_5821_0 : 3'h0;
  assign v_9019_0 = v_26_0 ? v_5807_0 : 3'h0;
  assign v_9020_0 = v_601_0 ? v_5800_0 : 3'h0;
  assign v_9021_0 = v_9022_0 | v_9023_0;
  assign v_9022_0 = v_607_0 ? v_5814_0 : 3'h0;
  assign v_9023_0 = v_26_0 ? v_5800_0 : 3'h0;
  assign v_9024_0 = v_601_0 ? v_5793_0 : 3'h0;
  assign v_9025_0 = v_9026_0 | v_9027_0;
  assign v_9026_0 = v_607_0 ? v_5807_0 : 3'h0;
  assign v_9027_0 = v_26_0 ? v_5793_0 : 3'h0;
  assign v_9028_0 = v_601_0 ? v_5786_0 : 3'h0;
  assign v_9029_0 = v_9030_0 | v_9031_0;
  assign v_9030_0 = v_607_0 ? v_5800_0 : 3'h0;
  assign v_9031_0 = v_26_0 ? v_5786_0 : 3'h0;
  assign v_9032_0 = v_601_0 ? v_5779_0 : 3'h0;
  assign v_9033_0 = v_9034_0 | v_9035_0;
  assign v_9034_0 = v_607_0 ? v_5793_0 : 3'h0;
  assign v_9035_0 = v_26_0 ? v_5779_0 : 3'h0;
  assign v_9036_0 = v_601_0 ? v_5772_0 : 3'h0;
  assign v_9037_0 = v_9038_0 | v_9039_0;
  assign v_9038_0 = v_607_0 ? v_5786_0 : 3'h0;
  assign v_9039_0 = v_26_0 ? v_5772_0 : 3'h0;
  assign v_9040_0 = v_601_0 ? v_5765_0 : 3'h0;
  assign v_9041_0 = v_9042_0 | v_9043_0;
  assign v_9042_0 = v_607_0 ? v_5779_0 : 3'h0;
  assign v_9043_0 = v_26_0 ? v_5765_0 : 3'h0;
  assign v_9044_0 = v_601_0 ? v_5758_0 : 3'h0;
  assign v_9045_0 = v_9046_0 | v_9047_0;
  assign v_9046_0 = v_607_0 ? v_5772_0 : 3'h0;
  assign v_9047_0 = v_26_0 ? v_5758_0 : 3'h0;
  assign v_9048_0 = v_601_0 ? v_5751_0 : 3'h0;
  assign v_9049_0 = v_9050_0 | v_9051_0;
  assign v_9050_0 = v_607_0 ? v_5765_0 : 3'h0;
  assign v_9051_0 = v_26_0 ? v_5751_0 : 3'h0;
  assign v_9052_0 = v_601_0 ? v_5744_0 : 3'h0;
  assign v_9053_0 = v_9054_0 | v_9055_0;
  assign v_9054_0 = v_607_0 ? v_5758_0 : 3'h0;
  assign v_9055_0 = v_26_0 ? v_5744_0 : 3'h0;
  assign v_9056_0 = v_601_0 ? v_5737_0 : 3'h0;
  assign v_9057_0 = v_9058_0 | v_9059_0;
  assign v_9058_0 = v_607_0 ? v_5751_0 : 3'h0;
  assign v_9059_0 = v_26_0 ? v_5737_0 : 3'h0;
  assign v_9060_0 = v_601_0 ? v_5730_0 : 3'h0;
  assign v_9061_0 = v_9062_0 | v_9063_0;
  assign v_9062_0 = v_607_0 ? v_5744_0 : 3'h0;
  assign v_9063_0 = v_26_0 ? v_5730_0 : 3'h0;
  assign v_9064_0 = v_601_0 ? v_5723_0 : 3'h0;
  assign v_9065_0 = v_9066_0 | v_9067_0;
  assign v_9066_0 = v_607_0 ? v_5737_0 : 3'h0;
  assign v_9067_0 = v_26_0 ? v_5723_0 : 3'h0;
  assign v_9068_0 = v_601_0 ? v_5716_0 : 3'h0;
  assign v_9069_0 = v_9070_0 | v_9071_0;
  assign v_9070_0 = v_607_0 ? v_5730_0 : 3'h0;
  assign v_9071_0 = v_26_0 ? v_5716_0 : 3'h0;
  assign v_9072_0 = v_601_0 ? v_5709_0 : 3'h0;
  assign v_9073_0 = v_9074_0 | v_9075_0;
  assign v_9074_0 = v_607_0 ? v_5723_0 : 3'h0;
  assign v_9075_0 = v_26_0 ? v_5709_0 : 3'h0;
  assign v_9076_0 = v_601_0 ? v_5702_0 : 3'h0;
  assign v_9077_0 = v_9078_0 | v_9079_0;
  assign v_9078_0 = v_607_0 ? v_5716_0 : 3'h0;
  assign v_9079_0 = v_26_0 ? v_5702_0 : 3'h0;
  assign v_9080_0 = v_601_0 ? v_5695_0 : 3'h0;
  assign v_9081_0 = v_9082_0 | v_9083_0;
  assign v_9082_0 = v_607_0 ? v_5709_0 : 3'h0;
  assign v_9083_0 = v_26_0 ? v_5695_0 : 3'h0;
  assign v_9084_0 = v_601_0 ? v_5688_0 : 3'h0;
  assign v_9085_0 = v_9086_0 | v_9087_0;
  assign v_9086_0 = v_607_0 ? v_5702_0 : 3'h0;
  assign v_9087_0 = v_26_0 ? v_5688_0 : 3'h0;
  assign v_9088_0 = v_601_0 ? v_5681_0 : 3'h0;
  assign v_9089_0 = v_9090_0 | v_9091_0;
  assign v_9090_0 = v_607_0 ? v_5695_0 : 3'h0;
  assign v_9091_0 = v_26_0 ? v_5681_0 : 3'h0;
  assign v_9092_0 = v_601_0 ? v_5674_0 : 3'h0;
  assign v_9093_0 = v_9094_0 | v_9095_0;
  assign v_9094_0 = v_607_0 ? v_5688_0 : 3'h0;
  assign v_9095_0 = v_26_0 ? v_5674_0 : 3'h0;
  assign v_9096_0 = v_601_0 ? v_5667_0 : 3'h0;
  assign v_9097_0 = v_9098_0 | v_9099_0;
  assign v_9098_0 = v_607_0 ? v_5681_0 : 3'h0;
  assign v_9099_0 = v_26_0 ? v_5667_0 : 3'h0;
  assign v_9100_0 = v_601_0 ? v_5660_0 : 3'h0;
  assign v_9101_0 = v_9102_0 | v_9103_0;
  assign v_9102_0 = v_607_0 ? v_5674_0 : 3'h0;
  assign v_9103_0 = v_26_0 ? v_5660_0 : 3'h0;
  assign v_9104_0 = v_601_0 ? v_5653_0 : 3'h0;
  assign v_9105_0 = v_9106_0 | v_9107_0;
  assign v_9106_0 = v_607_0 ? v_5667_0 : 3'h0;
  assign v_9107_0 = v_26_0 ? v_5653_0 : 3'h0;
  assign v_9108_0 = v_601_0 ? v_5646_0 : 3'h0;
  assign v_9109_0 = v_9110_0 | v_9111_0;
  assign v_9110_0 = v_607_0 ? v_5660_0 : 3'h0;
  assign v_9111_0 = v_26_0 ? v_5646_0 : 3'h0;
  assign v_9112_0 = v_601_0 ? v_5639_0 : 3'h0;
  assign v_9113_0 = v_9114_0 | v_9115_0;
  assign v_9114_0 = v_607_0 ? v_5653_0 : 3'h0;
  assign v_9115_0 = v_26_0 ? v_5639_0 : 3'h0;
  assign v_9116_0 = v_601_0 ? v_5632_0 : 3'h0;
  assign v_9117_0 = v_9118_0 | v_9119_0;
  assign v_9118_0 = v_607_0 ? v_5646_0 : 3'h0;
  assign v_9119_0 = v_26_0 ? v_5632_0 : 3'h0;
  assign v_9120_0 = v_601_0 ? v_5625_0 : 3'h0;
  assign v_9121_0 = v_9122_0 | v_9123_0;
  assign v_9122_0 = v_607_0 ? v_5639_0 : 3'h0;
  assign v_9123_0 = v_26_0 ? v_5625_0 : 3'h0;
  assign v_9124_0 = v_601_0 ? v_5618_0 : 3'h0;
  assign v_9125_0 = v_9126_0 | v_9127_0;
  assign v_9126_0 = v_607_0 ? v_5632_0 : 3'h0;
  assign v_9127_0 = v_26_0 ? v_5618_0 : 3'h0;
  assign v_9128_0 = v_601_0 ? v_5611_0 : 3'h0;
  assign v_9129_0 = v_9130_0 | v_9131_0;
  assign v_9130_0 = v_607_0 ? v_5625_0 : 3'h0;
  assign v_9131_0 = v_26_0 ? v_5611_0 : 3'h0;
  assign v_9132_0 = v_601_0 ? v_5604_0 : 3'h0;
  assign v_9133_0 = v_9134_0 | v_9135_0;
  assign v_9134_0 = v_607_0 ? v_5618_0 : 3'h0;
  assign v_9135_0 = v_26_0 ? v_5604_0 : 3'h0;
  assign v_9136_0 = v_601_0 ? v_5597_0 : 3'h0;
  assign v_9137_0 = v_9138_0 | v_9139_0;
  assign v_9138_0 = v_607_0 ? v_5611_0 : 3'h0;
  assign v_9139_0 = v_26_0 ? v_5597_0 : 3'h0;
  assign v_9140_0 = v_601_0 ? v_5590_0 : 3'h0;
  assign v_9141_0 = v_9142_0 | v_9143_0;
  assign v_9142_0 = v_607_0 ? v_5604_0 : 3'h0;
  assign v_9143_0 = v_26_0 ? v_5590_0 : 3'h0;
  assign v_9144_0 = v_601_0 ? v_5583_0 : 3'h0;
  assign v_9145_0 = v_9146_0 | v_9147_0;
  assign v_9146_0 = v_607_0 ? v_5597_0 : 3'h0;
  assign v_9147_0 = v_26_0 ? v_5583_0 : 3'h0;
  assign v_9148_0 = v_601_0 ? v_5576_0 : 3'h0;
  assign v_9149_0 = v_9150_0 | v_9151_0;
  assign v_9150_0 = v_607_0 ? v_5590_0 : 3'h0;
  assign v_9151_0 = v_26_0 ? v_5576_0 : 3'h0;
  assign v_9152_0 = v_601_0 ? v_5569_0 : 3'h0;
  assign v_9153_0 = v_9154_0 | v_9155_0;
  assign v_9154_0 = v_607_0 ? v_5583_0 : 3'h0;
  assign v_9155_0 = v_26_0 ? v_5569_0 : 3'h0;
  assign v_9156_0 = v_601_0 ? v_5562_0 : 3'h0;
  assign v_9157_0 = v_9158_0 | v_9159_0;
  assign v_9158_0 = v_607_0 ? v_5576_0 : 3'h0;
  assign v_9159_0 = v_26_0 ? v_5562_0 : 3'h0;
  assign v_9160_0 = v_601_0 ? v_5555_0 : 3'h0;
  assign v_9161_0 = v_9162_0 | v_9163_0;
  assign v_9162_0 = v_607_0 ? v_5569_0 : 3'h0;
  assign v_9163_0 = v_26_0 ? v_5555_0 : 3'h0;
  assign v_9164_0 = v_601_0 ? v_5548_0 : 3'h0;
  assign v_9165_0 = v_9166_0 | v_9167_0;
  assign v_9166_0 = v_607_0 ? v_5562_0 : 3'h0;
  assign v_9167_0 = v_26_0 ? v_5548_0 : 3'h0;
  assign v_9168_0 = v_601_0 ? v_5541_0 : 3'h0;
  assign v_9169_0 = v_9170_0 | v_9171_0;
  assign v_9170_0 = v_607_0 ? v_5555_0 : 3'h0;
  assign v_9171_0 = v_26_0 ? v_5541_0 : 3'h0;
  assign v_9172_0 = v_601_0 ? v_5534_0 : 3'h0;
  assign v_9173_0 = v_9174_0 | v_9175_0;
  assign v_9174_0 = v_607_0 ? v_5548_0 : 3'h0;
  assign v_9175_0 = v_26_0 ? v_5534_0 : 3'h0;
  assign v_9176_0 = v_601_0 ? v_5527_0 : 3'h0;
  assign v_9177_0 = v_9178_0 | v_9179_0;
  assign v_9178_0 = v_607_0 ? v_5541_0 : 3'h0;
  assign v_9179_0 = v_26_0 ? v_5527_0 : 3'h0;
  assign v_9180_0 = v_601_0 ? v_5520_0 : 3'h0;
  assign v_9181_0 = v_9182_0 | v_9183_0;
  assign v_9182_0 = v_607_0 ? v_5534_0 : 3'h0;
  assign v_9183_0 = v_26_0 ? v_5520_0 : 3'h0;
  assign v_9184_0 = v_601_0 ? v_5513_0 : 3'h0;
  assign v_9185_0 = v_9186_0 | v_9187_0;
  assign v_9186_0 = v_607_0 ? v_5527_0 : 3'h0;
  assign v_9187_0 = v_26_0 ? v_5513_0 : 3'h0;
  assign v_9188_0 = v_601_0 ? v_5506_0 : 3'h0;
  assign v_9189_0 = v_9190_0 | v_9191_0;
  assign v_9190_0 = v_607_0 ? v_5520_0 : 3'h0;
  assign v_9191_0 = v_26_0 ? v_5506_0 : 3'h0;
  assign v_9192_0 = v_601_0 ? v_5499_0 : 3'h0;
  assign v_9193_0 = v_9194_0 | v_9195_0;
  assign v_9194_0 = v_607_0 ? v_5513_0 : 3'h0;
  assign v_9195_0 = v_26_0 ? v_5499_0 : 3'h0;
  assign v_9196_0 = v_601_0 ? v_5492_0 : 3'h0;
  assign v_9197_0 = v_9198_0 | v_9199_0;
  assign v_9198_0 = v_607_0 ? v_5506_0 : 3'h0;
  assign v_9199_0 = v_26_0 ? v_5492_0 : 3'h0;
  assign v_9200_0 = v_601_0 ? v_5485_0 : 3'h0;
  assign v_9201_0 = v_9202_0 | v_9203_0;
  assign v_9202_0 = v_607_0 ? v_5499_0 : 3'h0;
  assign v_9203_0 = v_26_0 ? v_5485_0 : 3'h0;
  assign v_9204_0 = v_601_0 ? v_5478_0 : 3'h0;
  assign v_9205_0 = v_9206_0 | v_9207_0;
  assign v_9206_0 = v_607_0 ? v_5492_0 : 3'h0;
  assign v_9207_0 = v_26_0 ? v_5478_0 : 3'h0;
  assign v_9208_0 = v_601_0 ? v_5471_0 : 3'h0;
  assign v_9209_0 = v_9210_0 | v_9211_0;
  assign v_9210_0 = v_607_0 ? v_5485_0 : 3'h0;
  assign v_9211_0 = v_26_0 ? v_5471_0 : 3'h0;
  assign v_9212_0 = v_601_0 ? v_5464_0 : 3'h0;
  assign v_9213_0 = v_9214_0 | v_9215_0;
  assign v_9214_0 = v_607_0 ? v_5478_0 : 3'h0;
  assign v_9215_0 = v_26_0 ? v_5464_0 : 3'h0;
  assign v_9216_0 = v_601_0 ? v_5457_0 : 3'h0;
  assign v_9217_0 = v_9218_0 | v_9219_0;
  assign v_9218_0 = v_607_0 ? v_5471_0 : 3'h0;
  assign v_9219_0 = v_26_0 ? v_5457_0 : 3'h0;
  assign v_9220_0 = v_601_0 ? v_5450_0 : 3'h0;
  assign v_9221_0 = v_9222_0 | v_9223_0;
  assign v_9222_0 = v_607_0 ? v_5464_0 : 3'h0;
  assign v_9223_0 = v_26_0 ? v_5450_0 : 3'h0;
  assign v_9224_0 = v_601_0 ? v_5443_0 : 3'h0;
  assign v_9225_0 = v_9226_0 | v_9227_0;
  assign v_9226_0 = v_607_0 ? v_5457_0 : 3'h0;
  assign v_9227_0 = v_26_0 ? v_5443_0 : 3'h0;
  assign v_9228_0 = v_601_0 ? v_5436_0 : 3'h0;
  assign v_9229_0 = v_9230_0 | v_9231_0;
  assign v_9230_0 = v_607_0 ? v_5450_0 : 3'h0;
  assign v_9231_0 = v_26_0 ? v_5436_0 : 3'h0;
  assign v_9232_0 = v_601_0 ? v_5429_0 : 3'h0;
  assign v_9233_0 = v_9234_0 | v_9235_0;
  assign v_9234_0 = v_607_0 ? v_5443_0 : 3'h0;
  assign v_9235_0 = v_26_0 ? v_5429_0 : 3'h0;
  assign v_9236_0 = v_601_0 ? v_5422_0 : 3'h0;
  assign v_9237_0 = v_9238_0 | v_9239_0;
  assign v_9238_0 = v_607_0 ? v_5436_0 : 3'h0;
  assign v_9239_0 = v_26_0 ? v_5422_0 : 3'h0;
  assign v_9240_0 = v_601_0 ? v_5415_0 : 3'h0;
  assign v_9241_0 = v_9242_0 | v_9243_0;
  assign v_9242_0 = v_607_0 ? v_5429_0 : 3'h0;
  assign v_9243_0 = v_26_0 ? v_5415_0 : 3'h0;
  assign v_9244_0 = v_601_0 ? v_5408_0 : 3'h0;
  assign v_9245_0 = v_9246_0 | v_9247_0;
  assign v_9246_0 = v_607_0 ? v_5422_0 : 3'h0;
  assign v_9247_0 = v_26_0 ? v_5408_0 : 3'h0;
  assign v_9248_0 = v_601_0 ? v_5401_0 : 3'h0;
  assign v_9249_0 = v_9250_0 | v_9251_0;
  assign v_9250_0 = v_607_0 ? v_5415_0 : 3'h0;
  assign v_9251_0 = v_26_0 ? v_5401_0 : 3'h0;
  assign v_9252_0 = v_601_0 ? v_5394_0 : 3'h0;
  assign v_9253_0 = v_9254_0 | v_9255_0;
  assign v_9254_0 = v_607_0 ? v_5408_0 : 3'h0;
  assign v_9255_0 = v_26_0 ? v_5394_0 : 3'h0;
  assign v_9256_0 = v_601_0 ? v_5387_0 : 3'h0;
  assign v_9257_0 = v_9258_0 | v_9259_0;
  assign v_9258_0 = v_607_0 ? v_5401_0 : 3'h0;
  assign v_9259_0 = v_26_0 ? v_5387_0 : 3'h0;
  assign v_9260_0 = v_601_0 ? v_5380_0 : 3'h0;
  assign v_9261_0 = v_9262_0 | v_9263_0;
  assign v_9262_0 = v_607_0 ? v_5394_0 : 3'h0;
  assign v_9263_0 = v_26_0 ? v_5380_0 : 3'h0;
  assign v_9264_0 = v_601_0 ? v_5373_0 : 3'h0;
  assign v_9265_0 = v_9266_0 | v_9267_0;
  assign v_9266_0 = v_607_0 ? v_5387_0 : 3'h0;
  assign v_9267_0 = v_26_0 ? v_5373_0 : 3'h0;
  assign v_9268_0 = v_601_0 ? v_5366_0 : 3'h0;
  assign v_9269_0 = v_9270_0 | v_9271_0;
  assign v_9270_0 = v_607_0 ? v_5380_0 : 3'h0;
  assign v_9271_0 = v_26_0 ? v_5366_0 : 3'h0;
  assign v_9272_0 = v_601_0 ? v_5359_0 : 3'h0;
  assign v_9273_0 = v_9274_0 | v_9275_0;
  assign v_9274_0 = v_607_0 ? v_5373_0 : 3'h0;
  assign v_9275_0 = v_26_0 ? v_5359_0 : 3'h0;
  assign v_9276_0 = v_601_0 ? v_5352_0 : 3'h0;
  assign v_9277_0 = v_9278_0 | v_9279_0;
  assign v_9278_0 = v_607_0 ? v_5366_0 : 3'h0;
  assign v_9279_0 = v_26_0 ? v_5352_0 : 3'h0;
  assign v_9280_0 = v_601_0 ? v_5345_0 : 3'h0;
  assign v_9281_0 = v_9282_0 | v_9283_0;
  assign v_9282_0 = v_607_0 ? v_5359_0 : 3'h0;
  assign v_9283_0 = v_26_0 ? v_5345_0 : 3'h0;
  assign v_9284_0 = v_601_0 ? v_5338_0 : 3'h0;
  assign v_9285_0 = v_9286_0 | v_9287_0;
  assign v_9286_0 = v_607_0 ? v_5352_0 : 3'h0;
  assign v_9287_0 = v_26_0 ? v_5338_0 : 3'h0;
  assign v_9288_0 = v_601_0 ? v_5331_0 : 3'h0;
  assign v_9289_0 = v_9290_0 | v_9291_0;
  assign v_9290_0 = v_607_0 ? v_5345_0 : 3'h0;
  assign v_9291_0 = v_26_0 ? v_5331_0 : 3'h0;
  assign v_9292_0 = v_601_0 ? v_5324_0 : 3'h0;
  assign v_9293_0 = v_9294_0 | v_9295_0;
  assign v_9294_0 = v_607_0 ? v_5338_0 : 3'h0;
  assign v_9295_0 = v_26_0 ? v_5324_0 : 3'h0;
  assign v_9296_0 = v_601_0 ? v_5317_0 : 3'h0;
  assign v_9297_0 = v_9298_0 | v_9299_0;
  assign v_9298_0 = v_607_0 ? v_5331_0 : 3'h0;
  assign v_9299_0 = v_26_0 ? v_5317_0 : 3'h0;
  assign v_9300_0 = v_601_0 ? v_5310_0 : 3'h0;
  assign v_9301_0 = v_9302_0 | v_9303_0;
  assign v_9302_0 = v_607_0 ? v_5324_0 : 3'h0;
  assign v_9303_0 = v_26_0 ? v_5310_0 : 3'h0;
  assign v_9304_0 = v_601_0 ? v_5303_0 : 3'h0;
  assign v_9305_0 = v_9306_0 | v_9307_0;
  assign v_9306_0 = v_607_0 ? v_5317_0 : 3'h0;
  assign v_9307_0 = v_26_0 ? v_5303_0 : 3'h0;
  assign v_9308_0 = v_601_0 ? v_5296_0 : 3'h0;
  assign v_9309_0 = v_9310_0 | v_9311_0;
  assign v_9310_0 = v_607_0 ? v_5310_0 : 3'h0;
  assign v_9311_0 = v_26_0 ? v_5296_0 : 3'h0;
  assign v_9312_0 = v_601_0 ? v_5289_0 : 3'h0;
  assign v_9313_0 = v_9314_0 | v_9315_0;
  assign v_9314_0 = v_607_0 ? v_5303_0 : 3'h0;
  assign v_9315_0 = v_26_0 ? v_5289_0 : 3'h0;
  assign v_9316_0 = v_601_0 ? v_5282_0 : 3'h0;
  assign v_9317_0 = v_9318_0 | v_9319_0;
  assign v_9318_0 = v_607_0 ? v_5296_0 : 3'h0;
  assign v_9319_0 = v_26_0 ? v_5282_0 : 3'h0;
  assign v_9320_0 = v_601_0 ? v_5275_0 : 3'h0;
  assign v_9321_0 = v_9322_0 | v_9323_0;
  assign v_9322_0 = v_607_0 ? v_5289_0 : 3'h0;
  assign v_9323_0 = v_26_0 ? v_5275_0 : 3'h0;
  assign v_9324_0 = v_601_0 ? v_5268_0 : 3'h0;
  assign v_9325_0 = v_9326_0 | v_9327_0;
  assign v_9326_0 = v_607_0 ? v_5282_0 : 3'h0;
  assign v_9327_0 = v_26_0 ? v_5268_0 : 3'h0;
  assign v_9328_0 = v_601_0 ? v_5261_0 : 3'h0;
  assign v_9329_0 = v_9330_0 | v_9331_0;
  assign v_9330_0 = v_607_0 ? v_5275_0 : 3'h0;
  assign v_9331_0 = v_26_0 ? v_5261_0 : 3'h0;
  assign v_9332_0 = v_601_0 ? v_5254_0 : 3'h0;
  assign v_9333_0 = v_9334_0 | v_9335_0;
  assign v_9334_0 = v_607_0 ? v_5268_0 : 3'h0;
  assign v_9335_0 = v_26_0 ? v_5254_0 : 3'h0;
  assign v_9336_0 = v_601_0 ? v_5247_0 : 3'h0;
  assign v_9337_0 = v_9338_0 | v_9339_0;
  assign v_9338_0 = v_607_0 ? v_5261_0 : 3'h0;
  assign v_9339_0 = v_26_0 ? v_5247_0 : 3'h0;
  assign v_9340_0 = v_601_0 ? v_5240_0 : 3'h0;
  assign v_9341_0 = v_9342_0 | v_9343_0;
  assign v_9342_0 = v_607_0 ? v_5254_0 : 3'h0;
  assign v_9343_0 = v_26_0 ? v_5240_0 : 3'h0;
  assign v_9344_0 = v_601_0 ? v_5233_0 : 3'h0;
  assign v_9345_0 = v_9346_0 | v_9347_0;
  assign v_9346_0 = v_607_0 ? v_5247_0 : 3'h0;
  assign v_9347_0 = v_26_0 ? v_5233_0 : 3'h0;
  assign v_9348_0 = v_601_0 ? v_5226_0 : 3'h0;
  assign v_9349_0 = v_9350_0 | v_9351_0;
  assign v_9350_0 = v_607_0 ? v_5240_0 : 3'h0;
  assign v_9351_0 = v_26_0 ? v_5226_0 : 3'h0;
  assign v_9352_0 = v_601_0 ? v_5219_0 : 3'h0;
  assign v_9353_0 = v_9354_0 | v_9355_0;
  assign v_9354_0 = v_607_0 ? v_5233_0 : 3'h0;
  assign v_9355_0 = v_26_0 ? v_5219_0 : 3'h0;
  assign v_9356_0 = v_601_0 ? v_5212_0 : 3'h0;
  assign v_9357_0 = v_9358_0 | v_9359_0;
  assign v_9358_0 = v_607_0 ? v_5226_0 : 3'h0;
  assign v_9359_0 = v_26_0 ? v_5212_0 : 3'h0;
  assign v_9360_0 = v_601_0 ? v_5205_0 : 3'h0;
  assign v_9361_0 = v_9362_0 | v_9363_0;
  assign v_9362_0 = v_607_0 ? v_5219_0 : 3'h0;
  assign v_9363_0 = v_26_0 ? v_5205_0 : 3'h0;
  assign v_9364_0 = v_601_0 ? v_5198_0 : 3'h0;
  assign v_9365_0 = v_9366_0 | v_9367_0;
  assign v_9366_0 = v_607_0 ? v_5212_0 : 3'h0;
  assign v_9367_0 = v_26_0 ? v_5198_0 : 3'h0;
  assign v_9368_0 = v_601_0 ? v_5191_0 : 3'h0;
  assign v_9369_0 = v_9370_0 | v_9371_0;
  assign v_9370_0 = v_607_0 ? v_5205_0 : 3'h0;
  assign v_9371_0 = v_26_0 ? v_5191_0 : 3'h0;
  assign v_9372_0 = v_601_0 ? v_5184_0 : 3'h0;
  assign v_9373_0 = v_9374_0 | v_9375_0;
  assign v_9374_0 = v_607_0 ? v_5198_0 : 3'h0;
  assign v_9375_0 = v_26_0 ? v_5184_0 : 3'h0;
  assign v_9376_0 = v_601_0 ? v_5177_0 : 3'h0;
  assign v_9377_0 = v_9378_0 | v_9379_0;
  assign v_9378_0 = v_607_0 ? v_5191_0 : 3'h0;
  assign v_9379_0 = v_26_0 ? v_5177_0 : 3'h0;
  assign v_9380_0 = v_601_0 ? v_5170_0 : 3'h0;
  assign v_9381_0 = v_9382_0 | v_9383_0;
  assign v_9382_0 = v_607_0 ? v_5184_0 : 3'h0;
  assign v_9383_0 = v_26_0 ? v_5170_0 : 3'h0;
  assign v_9384_0 = v_601_0 ? v_5163_0 : 3'h0;
  assign v_9385_0 = v_9386_0 | v_9387_0;
  assign v_9386_0 = v_607_0 ? v_5177_0 : 3'h0;
  assign v_9387_0 = v_26_0 ? v_5163_0 : 3'h0;
  assign v_9388_0 = v_601_0 ? v_5156_0 : 3'h0;
  assign v_9389_0 = v_9390_0 | v_9391_0;
  assign v_9390_0 = v_607_0 ? v_5170_0 : 3'h0;
  assign v_9391_0 = v_26_0 ? v_5156_0 : 3'h0;
  assign v_9392_0 = v_601_0 ? v_5149_0 : 3'h0;
  assign v_9393_0 = v_9394_0 | v_9395_0;
  assign v_9394_0 = v_607_0 ? v_5163_0 : 3'h0;
  assign v_9395_0 = v_26_0 ? v_5149_0 : 3'h0;
  assign v_9396_0 = v_601_0 ? v_5142_0 : 3'h0;
  assign v_9397_0 = v_9398_0 | v_9399_0;
  assign v_9398_0 = v_607_0 ? v_5156_0 : 3'h0;
  assign v_9399_0 = v_26_0 ? v_5142_0 : 3'h0;
  assign v_9400_0 = v_601_0 ? v_5135_0 : 3'h0;
  assign v_9401_0 = v_9402_0 | v_9403_0;
  assign v_9402_0 = v_607_0 ? v_5149_0 : 3'h0;
  assign v_9403_0 = v_26_0 ? v_5135_0 : 3'h0;
  assign v_9404_0 = v_601_0 ? v_5128_0 : 3'h0;
  assign v_9405_0 = v_9406_0 | v_9407_0;
  assign v_9406_0 = v_607_0 ? v_5142_0 : 3'h0;
  assign v_9407_0 = v_26_0 ? v_5128_0 : 3'h0;
  assign v_9408_0 = v_601_0 ? v_5121_0 : 3'h0;
  assign v_9409_0 = v_9410_0 | v_9411_0;
  assign v_9410_0 = v_607_0 ? v_5135_0 : 3'h0;
  assign v_9411_0 = v_26_0 ? v_5121_0 : 3'h0;
  assign v_9412_0 = v_601_0 ? v_5114_0 : 3'h0;
  assign v_9413_0 = v_9414_0 | v_9415_0;
  assign v_9414_0 = v_607_0 ? v_5128_0 : 3'h0;
  assign v_9415_0 = v_26_0 ? v_5114_0 : 3'h0;
  assign v_9416_0 = v_601_0 ? v_5107_0 : 3'h0;
  assign v_9417_0 = v_9418_0 | v_9419_0;
  assign v_9418_0 = v_607_0 ? v_5121_0 : 3'h0;
  assign v_9419_0 = v_26_0 ? v_5107_0 : 3'h0;
  assign v_9420_0 = v_601_0 ? v_5100_0 : 3'h0;
  assign v_9421_0 = v_9422_0 | v_9423_0;
  assign v_9422_0 = v_607_0 ? v_5114_0 : 3'h0;
  assign v_9423_0 = v_26_0 ? v_5100_0 : 3'h0;
  assign v_9424_0 = v_601_0 ? v_5093_0 : 3'h0;
  assign v_9425_0 = v_9426_0 | v_9427_0;
  assign v_9426_0 = v_607_0 ? v_5107_0 : 3'h0;
  assign v_9427_0 = v_26_0 ? v_5093_0 : 3'h0;
  assign v_9428_0 = v_601_0 ? v_5086_0 : 3'h0;
  assign v_9429_0 = v_9430_0 | v_9431_0;
  assign v_9430_0 = v_607_0 ? v_5100_0 : 3'h0;
  assign v_9431_0 = v_26_0 ? v_5086_0 : 3'h0;
  assign v_9432_0 = v_601_0 ? v_5079_0 : 3'h0;
  assign v_9433_0 = v_9434_0 | v_9435_0;
  assign v_9434_0 = v_607_0 ? v_5093_0 : 3'h0;
  assign v_9435_0 = v_26_0 ? v_5079_0 : 3'h0;
  assign v_9436_0 = v_601_0 ? v_5072_0 : 3'h0;
  assign v_9437_0 = v_9438_0 | v_9439_0;
  assign v_9438_0 = v_607_0 ? v_5086_0 : 3'h0;
  assign v_9439_0 = v_26_0 ? v_5072_0 : 3'h0;
  assign v_9440_0 = v_601_0 ? v_5065_0 : 3'h0;
  assign v_9441_0 = v_9442_0 | v_9443_0;
  assign v_9442_0 = v_607_0 ? v_5079_0 : 3'h0;
  assign v_9443_0 = v_26_0 ? v_5065_0 : 3'h0;
  assign v_9444_0 = v_601_0 ? v_5058_0 : 3'h0;
  assign v_9445_0 = v_9446_0 | v_9447_0;
  assign v_9446_0 = v_607_0 ? v_5072_0 : 3'h0;
  assign v_9447_0 = v_26_0 ? v_5058_0 : 3'h0;
  assign v_9448_0 = v_601_0 ? v_5051_0 : 3'h0;
  assign v_9449_0 = v_9450_0 | v_9451_0;
  assign v_9450_0 = v_607_0 ? v_5065_0 : 3'h0;
  assign v_9451_0 = v_26_0 ? v_5051_0 : 3'h0;
  assign v_9452_0 = v_601_0 ? v_5044_0 : 3'h0;
  assign v_9453_0 = v_9454_0 | v_9455_0;
  assign v_9454_0 = v_607_0 ? v_5058_0 : 3'h0;
  assign v_9455_0 = v_26_0 ? v_5044_0 : 3'h0;
  assign v_9456_0 = v_601_0 ? v_5037_0 : 3'h0;
  assign v_9457_0 = v_9458_0 | v_9459_0;
  assign v_9458_0 = v_607_0 ? v_5051_0 : 3'h0;
  assign v_9459_0 = v_26_0 ? v_5037_0 : 3'h0;
  assign v_9460_0 = v_601_0 ? v_5030_0 : 3'h0;
  assign v_9461_0 = v_9462_0 | v_9463_0;
  assign v_9462_0 = v_607_0 ? v_5044_0 : 3'h0;
  assign v_9463_0 = v_26_0 ? v_5030_0 : 3'h0;
  assign v_9464_0 = v_601_0 ? v_5023_0 : 3'h0;
  assign v_9465_0 = v_9466_0 | v_9467_0;
  assign v_9466_0 = v_607_0 ? v_5037_0 : 3'h0;
  assign v_9467_0 = v_26_0 ? v_5023_0 : 3'h0;
  assign v_9468_0 = v_601_0 ? v_5016_0 : 3'h0;
  assign v_9469_0 = v_9470_0 | v_9471_0;
  assign v_9470_0 = v_607_0 ? v_5030_0 : 3'h0;
  assign v_9471_0 = v_26_0 ? v_5016_0 : 3'h0;
  assign v_9472_0 = v_601_0 ? v_5009_0 : 3'h0;
  assign v_9473_0 = v_9474_0 | v_9475_0;
  assign v_9474_0 = v_607_0 ? v_5023_0 : 3'h0;
  assign v_9475_0 = v_26_0 ? v_5009_0 : 3'h0;
  assign v_9476_0 = v_601_0 ? v_5002_0 : 3'h0;
  assign v_9477_0 = v_9478_0 | v_9479_0;
  assign v_9478_0 = v_607_0 ? v_5016_0 : 3'h0;
  assign v_9479_0 = v_26_0 ? v_5002_0 : 3'h0;
  assign v_9480_0 = v_601_0 ? v_4995_0 : 3'h0;
  assign v_9481_0 = v_9482_0 | v_9483_0;
  assign v_9482_0 = v_607_0 ? v_5009_0 : 3'h0;
  assign v_9483_0 = v_26_0 ? v_4995_0 : 3'h0;
  assign v_9484_0 = v_601_0 ? v_4988_0 : 3'h0;
  assign v_9485_0 = v_9486_0 | v_9487_0;
  assign v_9486_0 = v_607_0 ? v_5002_0 : 3'h0;
  assign v_9487_0 = v_26_0 ? v_4988_0 : 3'h0;
  assign v_9488_0 = v_601_0 ? v_4981_0 : 3'h0;
  assign v_9489_0 = v_9490_0 | v_9491_0;
  assign v_9490_0 = v_607_0 ? v_4995_0 : 3'h0;
  assign v_9491_0 = v_26_0 ? v_4981_0 : 3'h0;
  assign v_9492_0 = v_601_0 ? v_4974_0 : 3'h0;
  assign v_9493_0 = v_9494_0 | v_9495_0;
  assign v_9494_0 = v_607_0 ? v_4988_0 : 3'h0;
  assign v_9495_0 = v_26_0 ? v_4974_0 : 3'h0;
  assign v_9496_0 = v_601_0 ? v_4967_0 : 3'h0;
  assign v_9497_0 = v_9498_0 | v_9499_0;
  assign v_9498_0 = v_607_0 ? v_4981_0 : 3'h0;
  assign v_9499_0 = v_26_0 ? v_4967_0 : 3'h0;
  assign v_9500_0 = v_601_0 ? v_4960_0 : 3'h0;
  assign v_9501_0 = v_9502_0 | v_9503_0;
  assign v_9502_0 = v_607_0 ? v_4974_0 : 3'h0;
  assign v_9503_0 = v_26_0 ? v_4960_0 : 3'h0;
  assign v_9504_0 = v_601_0 ? v_4953_0 : 3'h0;
  assign v_9505_0 = v_9506_0 | v_9507_0;
  assign v_9506_0 = v_607_0 ? v_4967_0 : 3'h0;
  assign v_9507_0 = v_26_0 ? v_4953_0 : 3'h0;
  assign v_9508_0 = v_601_0 ? v_4946_0 : 3'h0;
  assign v_9509_0 = v_9510_0 | v_9511_0;
  assign v_9510_0 = v_607_0 ? v_4960_0 : 3'h0;
  assign v_9511_0 = v_26_0 ? v_4946_0 : 3'h0;
  assign v_9512_0 = v_601_0 ? v_4939_0 : 3'h0;
  assign v_9513_0 = v_9514_0 | v_9515_0;
  assign v_9514_0 = v_607_0 ? v_4953_0 : 3'h0;
  assign v_9515_0 = v_26_0 ? v_4939_0 : 3'h0;
  assign v_9516_0 = v_601_0 ? v_4932_0 : 3'h0;
  assign v_9517_0 = v_9518_0 | v_9519_0;
  assign v_9518_0 = v_607_0 ? v_4946_0 : 3'h0;
  assign v_9519_0 = v_26_0 ? v_4932_0 : 3'h0;
  assign v_9520_0 = v_601_0 ? v_4925_0 : 3'h0;
  assign v_9521_0 = v_9522_0 | v_9523_0;
  assign v_9522_0 = v_607_0 ? v_4939_0 : 3'h0;
  assign v_9523_0 = v_26_0 ? v_4925_0 : 3'h0;
  assign v_9524_0 = v_601_0 ? v_4918_0 : 3'h0;
  assign v_9525_0 = v_9526_0 | v_9527_0;
  assign v_9526_0 = v_607_0 ? v_4932_0 : 3'h0;
  assign v_9527_0 = v_26_0 ? v_4918_0 : 3'h0;
  assign v_9528_0 = v_601_0 ? v_4911_0 : 3'h0;
  assign v_9529_0 = v_9530_0 | v_9531_0;
  assign v_9530_0 = v_607_0 ? v_4925_0 : 3'h0;
  assign v_9531_0 = v_26_0 ? v_4911_0 : 3'h0;
  assign v_9532_0 = v_601_0 ? v_4904_0 : 3'h0;
  assign v_9533_0 = v_9534_0 | v_9535_0;
  assign v_9534_0 = v_607_0 ? v_4918_0 : 3'h0;
  assign v_9535_0 = v_26_0 ? v_4904_0 : 3'h0;
  assign v_9536_0 = v_601_0 ? v_4897_0 : 3'h0;
  assign v_9537_0 = v_9538_0 | v_9539_0;
  assign v_9538_0 = v_607_0 ? v_4911_0 : 3'h0;
  assign v_9539_0 = v_26_0 ? v_4897_0 : 3'h0;
  assign v_9540_0 = v_601_0 ? v_4890_0 : 3'h0;
  assign v_9541_0 = v_9542_0 | v_9543_0;
  assign v_9542_0 = v_607_0 ? v_4904_0 : 3'h0;
  assign v_9543_0 = v_26_0 ? v_4890_0 : 3'h0;
  assign v_9544_0 = v_601_0 ? v_4883_0 : 3'h0;
  assign v_9545_0 = v_9546_0 | v_9547_0;
  assign v_9546_0 = v_607_0 ? v_4897_0 : 3'h0;
  assign v_9547_0 = v_26_0 ? v_4883_0 : 3'h0;
  assign v_9548_0 = v_601_0 ? v_4876_0 : 3'h0;
  assign v_9549_0 = v_9550_0 | v_9551_0;
  assign v_9550_0 = v_607_0 ? v_4890_0 : 3'h0;
  assign v_9551_0 = v_26_0 ? v_4876_0 : 3'h0;
  assign v_9552_0 = v_601_0 ? v_4869_0 : 3'h0;
  assign v_9553_0 = v_9554_0 | v_9555_0;
  assign v_9554_0 = v_607_0 ? v_4883_0 : 3'h0;
  assign v_9555_0 = v_26_0 ? v_4869_0 : 3'h0;
  assign v_9556_0 = v_601_0 ? v_4862_0 : 3'h0;
  assign v_9557_0 = v_9558_0 | v_9559_0;
  assign v_9558_0 = v_607_0 ? v_4876_0 : 3'h0;
  assign v_9559_0 = v_26_0 ? v_4862_0 : 3'h0;
  assign v_9560_0 = v_601_0 ? v_4855_0 : 3'h0;
  assign v_9561_0 = v_9562_0 | v_9563_0;
  assign v_9562_0 = v_607_0 ? v_4869_0 : 3'h0;
  assign v_9563_0 = v_26_0 ? v_4855_0 : 3'h0;
  assign v_9564_0 = v_601_0 ? v_4848_0 : 3'h0;
  assign v_9565_0 = v_9566_0 | v_9567_0;
  assign v_9566_0 = v_607_0 ? v_4862_0 : 3'h0;
  assign v_9567_0 = v_26_0 ? v_4848_0 : 3'h0;
  assign v_9568_0 = v_601_0 ? v_4841_0 : 3'h0;
  assign v_9569_0 = v_9570_0 | v_9571_0;
  assign v_9570_0 = v_607_0 ? v_4855_0 : 3'h0;
  assign v_9571_0 = v_26_0 ? v_4841_0 : 3'h0;
  assign v_9572_0 = v_601_0 ? v_4834_0 : 3'h0;
  assign v_9573_0 = v_9574_0 | v_9575_0;
  assign v_9574_0 = v_607_0 ? v_4848_0 : 3'h0;
  assign v_9575_0 = v_26_0 ? v_4834_0 : 3'h0;
  assign v_9576_0 = v_601_0 ? v_4827_0 : 3'h0;
  assign v_9577_0 = v_9578_0 | v_9579_0;
  assign v_9578_0 = v_607_0 ? v_4841_0 : 3'h0;
  assign v_9579_0 = v_26_0 ? v_4827_0 : 3'h0;
  assign v_9580_0 = v_601_0 ? v_4820_0 : 3'h0;
  assign v_9581_0 = v_9582_0 | v_9583_0;
  assign v_9582_0 = v_607_0 ? v_4834_0 : 3'h0;
  assign v_9583_0 = v_26_0 ? v_4820_0 : 3'h0;
  assign v_9584_0 = v_601_0 ? v_4813_0 : 3'h0;
  assign v_9585_0 = v_9586_0 | v_9587_0;
  assign v_9586_0 = v_607_0 ? v_4827_0 : 3'h0;
  assign v_9587_0 = v_26_0 ? v_4813_0 : 3'h0;
  assign v_9588_0 = v_601_0 ? v_4806_0 : 3'h0;
  assign v_9589_0 = v_9590_0 | v_9591_0;
  assign v_9590_0 = v_607_0 ? v_4820_0 : 3'h0;
  assign v_9591_0 = v_26_0 ? v_4806_0 : 3'h0;
  assign v_9592_0 = v_601_0 ? v_4799_0 : 3'h0;
  assign v_9593_0 = v_9594_0 | v_9595_0;
  assign v_9594_0 = v_607_0 ? v_4813_0 : 3'h0;
  assign v_9595_0 = v_26_0 ? v_4799_0 : 3'h0;
  assign v_9596_0 = v_601_0 ? v_4792_0 : 3'h0;
  assign v_9597_0 = v_9598_0 | v_9599_0;
  assign v_9598_0 = v_607_0 ? v_4806_0 : 3'h0;
  assign v_9599_0 = v_26_0 ? v_4792_0 : 3'h0;
  assign v_9600_0 = v_601_0 ? v_4785_0 : 3'h0;
  assign v_9601_0 = v_9602_0 | v_9603_0;
  assign v_9602_0 = v_607_0 ? v_4799_0 : 3'h0;
  assign v_9603_0 = v_26_0 ? v_4785_0 : 3'h0;
  assign v_9604_0 = v_601_0 ? v_4778_0 : 3'h0;
  assign v_9605_0 = v_9606_0 | v_9607_0;
  assign v_9606_0 = v_607_0 ? v_4792_0 : 3'h0;
  assign v_9607_0 = v_26_0 ? v_4778_0 : 3'h0;
  assign v_9608_0 = v_601_0 ? v_4771_0 : 3'h0;
  assign v_9609_0 = v_9610_0 | v_9611_0;
  assign v_9610_0 = v_607_0 ? v_4785_0 : 3'h0;
  assign v_9611_0 = v_26_0 ? v_4771_0 : 3'h0;
  assign v_9612_0 = v_601_0 ? v_4764_0 : 3'h0;
  assign v_9613_0 = v_9614_0 | v_9615_0;
  assign v_9614_0 = v_607_0 ? v_4778_0 : 3'h0;
  assign v_9615_0 = v_26_0 ? v_4764_0 : 3'h0;
  assign v_9616_0 = v_601_0 ? v_4757_0 : 3'h0;
  assign v_9617_0 = v_9618_0 | v_9619_0;
  assign v_9618_0 = v_607_0 ? v_4771_0 : 3'h0;
  assign v_9619_0 = v_26_0 ? v_4757_0 : 3'h0;
  assign v_9620_0 = v_601_0 ? v_4750_0 : 3'h0;
  assign v_9621_0 = v_9622_0 | v_9623_0;
  assign v_9622_0 = v_607_0 ? v_4764_0 : 3'h0;
  assign v_9623_0 = v_26_0 ? v_4750_0 : 3'h0;
  assign v_9624_0 = v_601_0 ? v_4743_0 : 3'h0;
  assign v_9625_0 = v_9626_0 | v_9627_0;
  assign v_9626_0 = v_607_0 ? v_4757_0 : 3'h0;
  assign v_9627_0 = v_26_0 ? v_4743_0 : 3'h0;
  assign v_9628_0 = v_601_0 ? v_4736_0 : 3'h0;
  assign v_9629_0 = v_9630_0 | v_9631_0;
  assign v_9630_0 = v_607_0 ? v_4750_0 : 3'h0;
  assign v_9631_0 = v_26_0 ? v_4736_0 : 3'h0;
  assign v_9632_0 = v_601_0 ? v_4729_0 : 3'h0;
  assign v_9633_0 = v_9634_0 | v_9635_0;
  assign v_9634_0 = v_607_0 ? v_4743_0 : 3'h0;
  assign v_9635_0 = v_26_0 ? v_4729_0 : 3'h0;
  assign v_9636_0 = v_601_0 ? v_4722_0 : 3'h0;
  assign v_9637_0 = v_9638_0 | v_9639_0;
  assign v_9638_0 = v_607_0 ? v_4736_0 : 3'h0;
  assign v_9639_0 = v_26_0 ? v_4722_0 : 3'h0;
  assign v_9640_0 = v_601_0 ? v_4715_0 : 3'h0;
  assign v_9641_0 = v_9642_0 | v_9643_0;
  assign v_9642_0 = v_607_0 ? v_4729_0 : 3'h0;
  assign v_9643_0 = v_26_0 ? v_4715_0 : 3'h0;
  assign v_9644_0 = v_601_0 ? v_4708_0 : 3'h0;
  assign v_9645_0 = v_9646_0 | v_9647_0;
  assign v_9646_0 = v_607_0 ? v_4722_0 : 3'h0;
  assign v_9647_0 = v_26_0 ? v_4708_0 : 3'h0;
  assign v_9648_0 = v_601_0 ? v_4701_0 : 3'h0;
  assign v_9649_0 = v_9650_0 | v_9651_0;
  assign v_9650_0 = v_607_0 ? v_4715_0 : 3'h0;
  assign v_9651_0 = v_26_0 ? v_4701_0 : 3'h0;
  assign v_9652_0 = v_601_0 ? v_4694_0 : 3'h0;
  assign v_9653_0 = v_9654_0 | v_9655_0;
  assign v_9654_0 = v_607_0 ? v_4708_0 : 3'h0;
  assign v_9655_0 = v_26_0 ? v_4694_0 : 3'h0;
  assign v_9656_0 = v_601_0 ? v_4687_0 : 3'h0;
  assign v_9657_0 = v_9658_0 | v_9659_0;
  assign v_9658_0 = v_607_0 ? v_4701_0 : 3'h0;
  assign v_9659_0 = v_26_0 ? v_4687_0 : 3'h0;
  assign v_9660_0 = v_601_0 ? v_4680_0 : 3'h0;
  assign v_9661_0 = v_9662_0 | v_9663_0;
  assign v_9662_0 = v_607_0 ? v_4694_0 : 3'h0;
  assign v_9663_0 = v_26_0 ? v_4680_0 : 3'h0;
  assign v_9664_0 = v_601_0 ? v_4673_0 : 3'h0;
  assign v_9665_0 = v_9666_0 | v_9667_0;
  assign v_9666_0 = v_607_0 ? v_4687_0 : 3'h0;
  assign v_9667_0 = v_26_0 ? v_4673_0 : 3'h0;
  assign v_9668_0 = v_601_0 ? v_4666_0 : 3'h0;
  assign v_9669_0 = v_9670_0 | v_9671_0;
  assign v_9670_0 = v_607_0 ? v_4680_0 : 3'h0;
  assign v_9671_0 = v_26_0 ? v_4666_0 : 3'h0;
  assign v_9672_0 = v_601_0 ? v_4659_0 : 3'h0;
  assign v_9673_0 = v_9674_0 | v_9675_0;
  assign v_9674_0 = v_607_0 ? v_4673_0 : 3'h0;
  assign v_9675_0 = v_26_0 ? v_4659_0 : 3'h0;
  assign v_9676_0 = v_601_0 ? v_4652_0 : 3'h0;
  assign v_9677_0 = v_9678_0 | v_9679_0;
  assign v_9678_0 = v_607_0 ? v_4666_0 : 3'h0;
  assign v_9679_0 = v_26_0 ? v_4652_0 : 3'h0;
  assign v_9680_0 = v_601_0 ? v_4645_0 : 3'h0;
  assign v_9681_0 = v_9682_0 | v_9683_0;
  assign v_9682_0 = v_607_0 ? v_4659_0 : 3'h0;
  assign v_9683_0 = v_26_0 ? v_4645_0 : 3'h0;
  assign v_9684_0 = v_601_0 ? v_4638_0 : 3'h0;
  assign v_9685_0 = v_9686_0 | v_9687_0;
  assign v_9686_0 = v_607_0 ? v_4652_0 : 3'h0;
  assign v_9687_0 = v_26_0 ? v_4638_0 : 3'h0;
  assign v_9688_0 = v_601_0 ? v_4631_0 : 3'h0;
  assign v_9689_0 = v_9690_0 | v_9691_0;
  assign v_9690_0 = v_607_0 ? v_4645_0 : 3'h0;
  assign v_9691_0 = v_26_0 ? v_4631_0 : 3'h0;
  assign v_9692_0 = v_601_0 ? v_4624_0 : 3'h0;
  assign v_9693_0 = v_9694_0 | v_9695_0;
  assign v_9694_0 = v_607_0 ? v_4638_0 : 3'h0;
  assign v_9695_0 = v_26_0 ? v_4624_0 : 3'h0;
  assign v_9696_0 = v_601_0 ? v_4617_0 : 3'h0;
  assign v_9697_0 = v_9698_0 | v_9699_0;
  assign v_9698_0 = v_607_0 ? v_4631_0 : 3'h0;
  assign v_9699_0 = v_26_0 ? v_4617_0 : 3'h0;
  assign v_9700_0 = v_601_0 ? v_4610_0 : 3'h0;
  assign v_9701_0 = v_9702_0 | v_9703_0;
  assign v_9702_0 = v_607_0 ? v_4624_0 : 3'h0;
  assign v_9703_0 = v_26_0 ? v_4610_0 : 3'h0;
  assign v_9704_0 = v_601_0 ? v_4603_0 : 3'h0;
  assign v_9705_0 = v_9706_0 | v_9707_0;
  assign v_9706_0 = v_607_0 ? v_4617_0 : 3'h0;
  assign v_9707_0 = v_26_0 ? v_4603_0 : 3'h0;
  assign v_9708_0 = v_601_0 ? v_4596_0 : 3'h0;
  assign v_9709_0 = v_9710_0 | v_9711_0;
  assign v_9710_0 = v_607_0 ? v_4610_0 : 3'h0;
  assign v_9711_0 = v_26_0 ? v_4596_0 : 3'h0;
  assign v_9712_0 = v_601_0 ? v_4589_0 : 3'h0;
  assign v_9713_0 = v_9714_0 | v_9715_0;
  assign v_9714_0 = v_607_0 ? v_4603_0 : 3'h0;
  assign v_9715_0 = v_26_0 ? v_4589_0 : 3'h0;
  assign v_9716_0 = v_601_0 ? v_4582_0 : 3'h0;
  assign v_9717_0 = v_9718_0 | v_9719_0;
  assign v_9718_0 = v_607_0 ? v_4596_0 : 3'h0;
  assign v_9719_0 = v_26_0 ? v_4582_0 : 3'h0;
  assign v_9720_0 = v_601_0 ? v_4575_0 : 3'h0;
  assign v_9721_0 = v_9722_0 | v_9723_0;
  assign v_9722_0 = v_607_0 ? v_4589_0 : 3'h0;
  assign v_9723_0 = v_26_0 ? v_4575_0 : 3'h0;
  assign v_9724_0 = v_601_0 ? v_4568_0 : 3'h0;
  assign v_9725_0 = v_9726_0 | v_9727_0;
  assign v_9726_0 = v_607_0 ? v_4582_0 : 3'h0;
  assign v_9727_0 = v_26_0 ? v_4568_0 : 3'h0;
  assign v_9728_0 = v_601_0 ? v_4561_0 : 3'h0;
  assign v_9729_0 = v_9730_0 | v_9731_0;
  assign v_9730_0 = v_607_0 ? v_4575_0 : 3'h0;
  assign v_9731_0 = v_26_0 ? v_4561_0 : 3'h0;
  assign v_9732_0 = v_601_0 ? v_4554_0 : 3'h0;
  assign v_9733_0 = v_9734_0 | v_9735_0;
  assign v_9734_0 = v_607_0 ? v_4568_0 : 3'h0;
  assign v_9735_0 = v_26_0 ? v_4554_0 : 3'h0;
  assign v_9736_0 = v_601_0 ? v_4547_0 : 3'h0;
  assign v_9737_0 = v_9738_0 | v_9739_0;
  assign v_9738_0 = v_607_0 ? v_4561_0 : 3'h0;
  assign v_9739_0 = v_26_0 ? v_4547_0 : 3'h0;
  assign v_9740_0 = v_601_0 ? v_4540_0 : 3'h0;
  assign v_9741_0 = v_9742_0 | v_9743_0;
  assign v_9742_0 = v_607_0 ? v_4554_0 : 3'h0;
  assign v_9743_0 = v_26_0 ? v_4540_0 : 3'h0;
  assign v_9744_0 = v_601_0 ? v_4533_0 : 3'h0;
  assign v_9745_0 = v_9746_0 | v_9747_0;
  assign v_9746_0 = v_607_0 ? v_4547_0 : 3'h0;
  assign v_9747_0 = v_26_0 ? v_4533_0 : 3'h0;
  assign v_9748_0 = v_601_0 ? v_4526_0 : 3'h0;
  assign v_9749_0 = v_9750_0 | v_9751_0;
  assign v_9750_0 = v_607_0 ? v_4540_0 : 3'h0;
  assign v_9751_0 = v_26_0 ? v_4526_0 : 3'h0;
  assign v_9752_0 = v_601_0 ? v_4519_0 : 3'h0;
  assign v_9753_0 = v_9754_0 | v_9755_0;
  assign v_9754_0 = v_607_0 ? v_4533_0 : 3'h0;
  assign v_9755_0 = v_26_0 ? v_4519_0 : 3'h0;
  assign v_9756_0 = v_601_0 ? v_4512_0 : 3'h0;
  assign v_9757_0 = v_9758_0 | v_9759_0;
  assign v_9758_0 = v_607_0 ? v_4526_0 : 3'h0;
  assign v_9759_0 = v_26_0 ? v_4512_0 : 3'h0;
  assign v_9760_0 = v_601_0 ? v_4505_0 : 3'h0;
  assign v_9761_0 = v_9762_0 | v_9763_0;
  assign v_9762_0 = v_607_0 ? v_4519_0 : 3'h0;
  assign v_9763_0 = v_26_0 ? v_4505_0 : 3'h0;
  assign v_9764_0 = v_601_0 ? v_4498_0 : 3'h0;
  assign v_9765_0 = v_9766_0 | v_9767_0;
  assign v_9766_0 = v_607_0 ? v_4512_0 : 3'h0;
  assign v_9767_0 = v_26_0 ? v_4498_0 : 3'h0;
  assign v_9768_0 = v_601_0 ? v_4491_0 : 3'h0;
  assign v_9769_0 = v_9770_0 | v_9771_0;
  assign v_9770_0 = v_607_0 ? v_4505_0 : 3'h0;
  assign v_9771_0 = v_26_0 ? v_4491_0 : 3'h0;
  assign v_9772_0 = v_601_0 ? v_4484_0 : 3'h0;
  assign v_9773_0 = v_9774_0 | v_9775_0;
  assign v_9774_0 = v_607_0 ? v_4498_0 : 3'h0;
  assign v_9775_0 = v_26_0 ? v_4484_0 : 3'h0;
  assign v_9776_0 = v_601_0 ? v_4477_0 : 3'h0;
  assign v_9777_0 = v_9778_0 | v_9779_0;
  assign v_9778_0 = v_607_0 ? v_4491_0 : 3'h0;
  assign v_9779_0 = v_26_0 ? v_4477_0 : 3'h0;
  assign v_9780_0 = v_601_0 ? v_4470_0 : 3'h0;
  assign v_9781_0 = v_9782_0 | v_9783_0;
  assign v_9782_0 = v_607_0 ? v_4484_0 : 3'h0;
  assign v_9783_0 = v_26_0 ? v_4470_0 : 3'h0;
  assign v_9784_0 = v_601_0 ? v_4463_0 : 3'h0;
  assign v_9785_0 = v_9786_0 | v_9787_0;
  assign v_9786_0 = v_607_0 ? v_4477_0 : 3'h0;
  assign v_9787_0 = v_26_0 ? v_4463_0 : 3'h0;
  assign v_9788_0 = v_601_0 ? v_4456_0 : 3'h0;
  assign v_9789_0 = v_9790_0 | v_9791_0;
  assign v_9790_0 = v_607_0 ? v_4470_0 : 3'h0;
  assign v_9791_0 = v_26_0 ? v_4456_0 : 3'h0;
  assign v_9792_0 = v_601_0 ? v_4449_0 : 3'h0;
  assign v_9793_0 = v_9794_0 | v_9795_0;
  assign v_9794_0 = v_607_0 ? v_4463_0 : 3'h0;
  assign v_9795_0 = v_26_0 ? v_4449_0 : 3'h0;
  assign v_9796_0 = v_601_0 ? v_4442_0 : 3'h0;
  assign v_9797_0 = v_9798_0 | v_9799_0;
  assign v_9798_0 = v_607_0 ? v_4456_0 : 3'h0;
  assign v_9799_0 = v_26_0 ? v_4442_0 : 3'h0;
  assign v_9800_0 = v_601_0 ? v_4435_0 : 3'h0;
  assign v_9801_0 = v_9802_0 | v_9803_0;
  assign v_9802_0 = v_607_0 ? v_4449_0 : 3'h0;
  assign v_9803_0 = v_26_0 ? v_4435_0 : 3'h0;
  assign v_9804_0 = v_601_0 ? v_4428_0 : 3'h0;
  assign v_9805_0 = v_9806_0 | v_9807_0;
  assign v_9806_0 = v_607_0 ? v_4442_0 : 3'h0;
  assign v_9807_0 = v_26_0 ? v_4428_0 : 3'h0;
  assign v_9808_0 = v_601_0 ? v_4421_0 : 3'h0;
  assign v_9809_0 = v_9810_0 | v_9811_0;
  assign v_9810_0 = v_607_0 ? v_4435_0 : 3'h0;
  assign v_9811_0 = v_26_0 ? v_4421_0 : 3'h0;
  assign v_9812_0 = v_601_0 ? v_4414_0 : 3'h0;
  assign v_9813_0 = v_9814_0 | v_9815_0;
  assign v_9814_0 = v_607_0 ? v_4428_0 : 3'h0;
  assign v_9815_0 = v_26_0 ? v_4414_0 : 3'h0;
  assign v_9816_0 = v_601_0 ? v_4407_0 : 3'h0;
  assign v_9817_0 = v_9818_0 | v_9819_0;
  assign v_9818_0 = v_607_0 ? v_4421_0 : 3'h0;
  assign v_9819_0 = v_26_0 ? v_4407_0 : 3'h0;
  assign v_9820_0 = v_601_0 ? v_4400_0 : 3'h0;
  assign v_9821_0 = v_9822_0 | v_9823_0;
  assign v_9822_0 = v_607_0 ? v_4414_0 : 3'h0;
  assign v_9823_0 = v_26_0 ? v_4400_0 : 3'h0;
  assign v_9824_0 = v_601_0 ? v_4393_0 : 3'h0;
  assign v_9825_0 = v_9826_0 | v_9827_0;
  assign v_9826_0 = v_607_0 ? v_4407_0 : 3'h0;
  assign v_9827_0 = v_26_0 ? v_4393_0 : 3'h0;
  assign v_9828_0 = v_601_0 ? v_4386_0 : 3'h0;
  assign v_9829_0 = v_9830_0 | v_9831_0;
  assign v_9830_0 = v_607_0 ? v_4400_0 : 3'h0;
  assign v_9831_0 = v_26_0 ? v_4386_0 : 3'h0;
  assign v_9832_0 = v_601_0 ? v_4379_0 : 3'h0;
  assign v_9833_0 = v_9834_0 | v_9835_0;
  assign v_9834_0 = v_607_0 ? v_4393_0 : 3'h0;
  assign v_9835_0 = v_26_0 ? v_4379_0 : 3'h0;
  assign v_9836_0 = v_601_0 ? v_4372_0 : 3'h0;
  assign v_9837_0 = v_9838_0 | v_9839_0;
  assign v_9838_0 = v_607_0 ? v_4386_0 : 3'h0;
  assign v_9839_0 = v_26_0 ? v_4372_0 : 3'h0;
  assign v_9840_0 = v_601_0 ? v_4365_0 : 3'h0;
  assign v_9841_0 = v_9842_0 | v_9843_0;
  assign v_9842_0 = v_607_0 ? v_4379_0 : 3'h0;
  assign v_9843_0 = v_26_0 ? v_4365_0 : 3'h0;
  assign v_9844_0 = v_601_0 ? v_4358_0 : 3'h0;
  assign v_9845_0 = v_9846_0 | v_9847_0;
  assign v_9846_0 = v_607_0 ? v_4372_0 : 3'h0;
  assign v_9847_0 = v_26_0 ? v_4358_0 : 3'h0;
  assign v_9848_0 = v_601_0 ? v_4351_0 : 3'h0;
  assign v_9849_0 = v_9850_0 | v_9851_0;
  assign v_9850_0 = v_607_0 ? v_4365_0 : 3'h0;
  assign v_9851_0 = v_26_0 ? v_4351_0 : 3'h0;
  assign v_9852_0 = v_601_0 ? v_4344_0 : 3'h0;
  assign v_9853_0 = v_9854_0 | v_9855_0;
  assign v_9854_0 = v_607_0 ? v_4358_0 : 3'h0;
  assign v_9855_0 = v_26_0 ? v_4344_0 : 3'h0;
  assign v_9856_0 = v_601_0 ? v_4337_0 : 3'h0;
  assign v_9857_0 = v_9858_0 | v_9859_0;
  assign v_9858_0 = v_607_0 ? v_4351_0 : 3'h0;
  assign v_9859_0 = v_26_0 ? v_4337_0 : 3'h0;
  assign v_9860_0 = v_601_0 ? v_4330_0 : 3'h0;
  assign v_9861_0 = v_9862_0 | v_9863_0;
  assign v_9862_0 = v_607_0 ? v_4344_0 : 3'h0;
  assign v_9863_0 = v_26_0 ? v_4330_0 : 3'h0;
  assign v_9864_0 = v_601_0 ? v_4323_0 : 3'h0;
  assign v_9865_0 = v_9866_0 | v_9867_0;
  assign v_9866_0 = v_607_0 ? v_4337_0 : 3'h0;
  assign v_9867_0 = v_26_0 ? v_4323_0 : 3'h0;
  assign v_9868_0 = v_601_0 ? v_4316_0 : 3'h0;
  assign v_9869_0 = v_9870_0 | v_9871_0;
  assign v_9870_0 = v_607_0 ? v_4330_0 : 3'h0;
  assign v_9871_0 = v_26_0 ? v_4316_0 : 3'h0;
  assign v_9872_0 = v_601_0 ? v_4309_0 : 3'h0;
  assign v_9873_0 = v_9874_0 | v_9875_0;
  assign v_9874_0 = v_607_0 ? v_4323_0 : 3'h0;
  assign v_9875_0 = v_26_0 ? v_4309_0 : 3'h0;
  assign v_9876_0 = v_601_0 ? v_4302_0 : 3'h0;
  assign v_9877_0 = v_9878_0 | v_9879_0;
  assign v_9878_0 = v_607_0 ? v_4316_0 : 3'h0;
  assign v_9879_0 = v_26_0 ? v_4302_0 : 3'h0;
  assign v_9880_0 = v_601_0 ? v_4295_0 : 3'h0;
  assign v_9881_0 = v_9882_0 | v_9883_0;
  assign v_9882_0 = v_607_0 ? v_4309_0 : 3'h0;
  assign v_9883_0 = v_26_0 ? v_4295_0 : 3'h0;
  assign v_9884_0 = v_601_0 ? v_4288_0 : 3'h0;
  assign v_9885_0 = v_9886_0 | v_9887_0;
  assign v_9886_0 = v_607_0 ? v_4302_0 : 3'h0;
  assign v_9887_0 = v_26_0 ? v_4288_0 : 3'h0;
  assign v_9888_0 = v_601_0 ? v_4281_0 : 3'h0;
  assign v_9889_0 = v_9890_0 | v_9891_0;
  assign v_9890_0 = v_607_0 ? v_4295_0 : 3'h0;
  assign v_9891_0 = v_26_0 ? v_4281_0 : 3'h0;
  assign v_9892_0 = v_601_0 ? v_4274_0 : 3'h0;
  assign v_9893_0 = v_9894_0 | v_9895_0;
  assign v_9894_0 = v_607_0 ? v_4288_0 : 3'h0;
  assign v_9895_0 = v_26_0 ? v_4274_0 : 3'h0;
  assign v_9896_0 = v_601_0 ? v_4267_0 : 3'h0;
  assign v_9897_0 = v_9898_0 | v_9899_0;
  assign v_9898_0 = v_607_0 ? v_4281_0 : 3'h0;
  assign v_9899_0 = v_26_0 ? v_4267_0 : 3'h0;
  assign v_9900_0 = v_601_0 ? v_4260_0 : 3'h0;
  assign v_9901_0 = v_9902_0 | v_9903_0;
  assign v_9902_0 = v_607_0 ? v_4274_0 : 3'h0;
  assign v_9903_0 = v_26_0 ? v_4260_0 : 3'h0;
  assign v_9904_0 = v_601_0 ? v_4253_0 : 3'h0;
  assign v_9905_0 = v_9906_0 | v_9907_0;
  assign v_9906_0 = v_607_0 ? v_4267_0 : 3'h0;
  assign v_9907_0 = v_26_0 ? v_4253_0 : 3'h0;
  assign v_9908_0 = v_601_0 ? v_4246_0 : 3'h0;
  assign v_9909_0 = v_9910_0 | v_9911_0;
  assign v_9910_0 = v_607_0 ? v_4260_0 : 3'h0;
  assign v_9911_0 = v_26_0 ? v_4246_0 : 3'h0;
  assign v_9912_0 = v_601_0 ? v_4239_0 : 3'h0;
  assign v_9913_0 = v_9914_0 | v_9915_0;
  assign v_9914_0 = v_607_0 ? v_4253_0 : 3'h0;
  assign v_9915_0 = v_26_0 ? v_4239_0 : 3'h0;
  assign v_9916_0 = v_601_0 ? v_4232_0 : 3'h0;
  assign v_9917_0 = v_9918_0 | v_9919_0;
  assign v_9918_0 = v_607_0 ? v_4246_0 : 3'h0;
  assign v_9919_0 = v_26_0 ? v_4232_0 : 3'h0;
  assign v_9920_0 = v_601_0 ? v_4225_0 : 3'h0;
  assign v_9921_0 = v_9922_0 | v_9923_0;
  assign v_9922_0 = v_607_0 ? v_4239_0 : 3'h0;
  assign v_9923_0 = v_26_0 ? v_4225_0 : 3'h0;
  assign v_9924_0 = v_601_0 ? v_4218_0 : 3'h0;
  assign v_9925_0 = v_9926_0 | v_9927_0;
  assign v_9926_0 = v_607_0 ? v_4232_0 : 3'h0;
  assign v_9927_0 = v_26_0 ? v_4218_0 : 3'h0;
  assign v_9928_0 = v_601_0 ? v_4211_0 : 3'h0;
  assign v_9929_0 = v_9930_0 | v_9931_0;
  assign v_9930_0 = v_607_0 ? v_4225_0 : 3'h0;
  assign v_9931_0 = v_26_0 ? v_4211_0 : 3'h0;
  assign v_9932_0 = v_601_0 ? v_4204_0 : 3'h0;
  assign v_9933_0 = v_9934_0 | v_9935_0;
  assign v_9934_0 = v_607_0 ? v_4218_0 : 3'h0;
  assign v_9935_0 = v_26_0 ? v_4204_0 : 3'h0;
  assign v_9936_0 = v_601_0 ? v_4197_0 : 3'h0;
  assign v_9937_0 = v_9938_0 | v_9939_0;
  assign v_9938_0 = v_607_0 ? v_4211_0 : 3'h0;
  assign v_9939_0 = v_26_0 ? v_4197_0 : 3'h0;
  assign v_9940_0 = v_601_0 ? v_4190_0 : 3'h0;
  assign v_9941_0 = v_9942_0 | v_9943_0;
  assign v_9942_0 = v_607_0 ? v_4204_0 : 3'h0;
  assign v_9943_0 = v_26_0 ? v_4190_0 : 3'h0;
  assign v_9944_0 = v_601_0 ? v_4183_0 : 3'h0;
  assign v_9945_0 = v_9946_0 | v_9947_0;
  assign v_9946_0 = v_607_0 ? v_4197_0 : 3'h0;
  assign v_9947_0 = v_26_0 ? v_4183_0 : 3'h0;
  assign v_9948_0 = v_601_0 ? v_4176_0 : 3'h0;
  assign v_9949_0 = v_9950_0 | v_9951_0;
  assign v_9950_0 = v_607_0 ? v_4190_0 : 3'h0;
  assign v_9951_0 = v_26_0 ? v_4176_0 : 3'h0;
  assign v_9952_0 = v_601_0 ? v_4169_0 : 3'h0;
  assign v_9953_0 = v_9954_0 | v_9955_0;
  assign v_9954_0 = v_607_0 ? v_4183_0 : 3'h0;
  assign v_9955_0 = v_26_0 ? v_4169_0 : 3'h0;
  assign v_9956_0 = v_601_0 ? v_4162_0 : 3'h0;
  assign v_9957_0 = v_9958_0 | v_9959_0;
  assign v_9958_0 = v_607_0 ? v_4176_0 : 3'h0;
  assign v_9959_0 = v_26_0 ? v_4162_0 : 3'h0;
  assign v_9960_0 = v_601_0 ? v_4155_0 : 3'h0;
  assign v_9961_0 = v_9962_0 | v_9963_0;
  assign v_9962_0 = v_607_0 ? v_4169_0 : 3'h0;
  assign v_9963_0 = v_26_0 ? v_4155_0 : 3'h0;
  assign v_9964_0 = v_601_0 ? v_4148_0 : 3'h0;
  assign v_9965_0 = v_9966_0 | v_9967_0;
  assign v_9966_0 = v_607_0 ? v_4162_0 : 3'h0;
  assign v_9967_0 = v_26_0 ? v_4148_0 : 3'h0;
  assign v_9968_0 = v_601_0 ? v_4141_0 : 3'h0;
  assign v_9969_0 = v_9970_0 | v_9971_0;
  assign v_9970_0 = v_607_0 ? v_4155_0 : 3'h0;
  assign v_9971_0 = v_26_0 ? v_4141_0 : 3'h0;
  assign v_9972_0 = v_601_0 ? v_4134_0 : 3'h0;
  assign v_9973_0 = v_9974_0 | v_9975_0;
  assign v_9974_0 = v_607_0 ? v_4148_0 : 3'h0;
  assign v_9975_0 = v_26_0 ? v_4134_0 : 3'h0;
  assign v_9976_0 = v_601_0 ? v_4127_0 : 3'h0;
  assign v_9977_0 = v_9978_0 | v_9979_0;
  assign v_9978_0 = v_607_0 ? v_4141_0 : 3'h0;
  assign v_9979_0 = v_26_0 ? v_4127_0 : 3'h0;
  assign v_9980_0 = v_601_0 ? v_4120_0 : 3'h0;
  assign v_9981_0 = v_9982_0 | v_9983_0;
  assign v_9982_0 = v_607_0 ? v_4134_0 : 3'h0;
  assign v_9983_0 = v_26_0 ? v_4120_0 : 3'h0;
  assign v_9984_0 = v_601_0 ? v_4113_0 : 3'h0;
  assign v_9985_0 = v_9986_0 | v_9987_0;
  assign v_9986_0 = v_607_0 ? v_4127_0 : 3'h0;
  assign v_9987_0 = v_26_0 ? v_4113_0 : 3'h0;
  assign v_9988_0 = v_601_0 ? v_4106_0 : 3'h0;
  assign v_9989_0 = v_9990_0 | v_9991_0;
  assign v_9990_0 = v_607_0 ? v_4120_0 : 3'h0;
  assign v_9991_0 = v_26_0 ? v_4106_0 : 3'h0;
  assign v_9992_0 = v_601_0 ? v_4099_0 : 3'h0;
  assign v_9993_0 = v_9994_0 | v_9995_0;
  assign v_9994_0 = v_607_0 ? v_4113_0 : 3'h0;
  assign v_9995_0 = v_26_0 ? v_4099_0 : 3'h0;
  assign v_9996_0 = v_601_0 ? v_4092_0 : 3'h0;
  assign v_9997_0 = v_9998_0 | v_9999_0;
  assign v_9998_0 = v_607_0 ? v_4106_0 : 3'h0;
  assign v_9999_0 = v_26_0 ? v_4092_0 : 3'h0;
  assign v_10000_0 = v_601_0 ? v_4085_0 : 3'h0;
  assign v_10001_0 = v_10002_0 | v_10003_0;
  assign v_10002_0 = v_607_0 ? v_4099_0 : 3'h0;
  assign v_10003_0 = v_26_0 ? v_4085_0 : 3'h0;
  assign v_10004_0 = v_601_0 ? v_4078_0 : 3'h0;
  assign v_10005_0 = v_10006_0 | v_10007_0;
  assign v_10006_0 = v_607_0 ? v_4092_0 : 3'h0;
  assign v_10007_0 = v_26_0 ? v_4078_0 : 3'h0;
  assign v_10008_0 = v_601_0 ? v_4071_0 : 3'h0;
  assign v_10009_0 = v_10010_0 | v_10011_0;
  assign v_10010_0 = v_607_0 ? v_4085_0 : 3'h0;
  assign v_10011_0 = v_26_0 ? v_4071_0 : 3'h0;
  assign v_10012_0 = v_601_0 ? v_4064_0 : 3'h0;
  assign v_10013_0 = v_10014_0 | v_10015_0;
  assign v_10014_0 = v_607_0 ? v_4078_0 : 3'h0;
  assign v_10015_0 = v_26_0 ? v_4064_0 : 3'h0;
  assign v_10016_0 = v_601_0 ? v_4057_0 : 3'h0;
  assign v_10017_0 = v_10018_0 | v_10019_0;
  assign v_10018_0 = v_607_0 ? v_4071_0 : 3'h0;
  assign v_10019_0 = v_26_0 ? v_4057_0 : 3'h0;
  assign v_10020_0 = v_601_0 ? v_4050_0 : 3'h0;
  assign v_10021_0 = v_10022_0 | v_10023_0;
  assign v_10022_0 = v_607_0 ? v_4064_0 : 3'h0;
  assign v_10023_0 = v_26_0 ? v_4050_0 : 3'h0;
  assign v_10024_0 = v_601_0 ? v_4043_0 : 3'h0;
  assign v_10025_0 = v_10026_0 | v_10027_0;
  assign v_10026_0 = v_607_0 ? v_4057_0 : 3'h0;
  assign v_10027_0 = v_26_0 ? v_4043_0 : 3'h0;
  assign v_10028_0 = v_601_0 ? v_4036_0 : 3'h0;
  assign v_10029_0 = v_10030_0 | v_10031_0;
  assign v_10030_0 = v_607_0 ? v_4050_0 : 3'h0;
  assign v_10031_0 = v_26_0 ? v_4036_0 : 3'h0;
  assign v_10032_0 = v_601_0 ? v_4029_0 : 3'h0;
  assign v_10033_0 = v_10034_0 | v_10035_0;
  assign v_10034_0 = v_607_0 ? v_4043_0 : 3'h0;
  assign v_10035_0 = v_26_0 ? v_4029_0 : 3'h0;
  assign v_10036_0 = v_601_0 ? v_4022_0 : 3'h0;
  assign v_10037_0 = v_10038_0 | v_10039_0;
  assign v_10038_0 = v_607_0 ? v_4036_0 : 3'h0;
  assign v_10039_0 = v_26_0 ? v_4022_0 : 3'h0;
  assign v_10040_0 = v_601_0 ? v_4015_0 : 3'h0;
  assign v_10041_0 = v_10042_0 | v_10043_0;
  assign v_10042_0 = v_607_0 ? v_4029_0 : 3'h0;
  assign v_10043_0 = v_26_0 ? v_4015_0 : 3'h0;
  assign v_10044_0 = v_601_0 ? v_4008_0 : 3'h0;
  assign v_10045_0 = v_10046_0 | v_10047_0;
  assign v_10046_0 = v_607_0 ? v_4022_0 : 3'h0;
  assign v_10047_0 = v_26_0 ? v_4008_0 : 3'h0;
  assign v_10048_0 = v_601_0 ? v_4001_0 : 3'h0;
  assign v_10049_0 = v_10050_0 | v_10051_0;
  assign v_10050_0 = v_607_0 ? v_4015_0 : 3'h0;
  assign v_10051_0 = v_26_0 ? v_4001_0 : 3'h0;
  assign v_10052_0 = v_601_0 ? v_3994_0 : 3'h0;
  assign v_10053_0 = v_10054_0 | v_10055_0;
  assign v_10054_0 = v_607_0 ? v_4008_0 : 3'h0;
  assign v_10055_0 = v_26_0 ? v_3994_0 : 3'h0;
  assign v_10056_0 = v_601_0 ? v_3987_0 : 3'h0;
  assign v_10057_0 = v_10058_0 | v_10059_0;
  assign v_10058_0 = v_607_0 ? v_4001_0 : 3'h0;
  assign v_10059_0 = v_26_0 ? v_3987_0 : 3'h0;
  assign v_10060_0 = v_601_0 ? v_3980_0 : 3'h0;
  assign v_10061_0 = v_10062_0 | v_10063_0;
  assign v_10062_0 = v_607_0 ? v_3994_0 : 3'h0;
  assign v_10063_0 = v_26_0 ? v_3980_0 : 3'h0;
  assign v_10064_0 = v_601_0 ? v_3973_0 : 3'h0;
  assign v_10065_0 = v_10066_0 | v_10067_0;
  assign v_10066_0 = v_607_0 ? v_3987_0 : 3'h0;
  assign v_10067_0 = v_26_0 ? v_3973_0 : 3'h0;
  assign v_10068_0 = v_601_0 ? v_3966_0 : 3'h0;
  assign v_10069_0 = v_10070_0 | v_10071_0;
  assign v_10070_0 = v_607_0 ? v_3980_0 : 3'h0;
  assign v_10071_0 = v_26_0 ? v_3966_0 : 3'h0;
  assign v_10072_0 = v_601_0 ? v_3959_0 : 3'h0;
  assign v_10073_0 = v_10074_0 | v_10075_0;
  assign v_10074_0 = v_607_0 ? v_3973_0 : 3'h0;
  assign v_10075_0 = v_26_0 ? v_3959_0 : 3'h0;
  assign v_10076_0 = v_601_0 ? v_3952_0 : 3'h0;
  assign v_10077_0 = v_10078_0 | v_10079_0;
  assign v_10078_0 = v_607_0 ? v_3966_0 : 3'h0;
  assign v_10079_0 = v_26_0 ? v_3952_0 : 3'h0;
  assign v_10080_0 = v_601_0 ? v_3945_0 : 3'h0;
  assign v_10081_0 = v_10082_0 | v_10083_0;
  assign v_10082_0 = v_607_0 ? v_3959_0 : 3'h0;
  assign v_10083_0 = v_26_0 ? v_3945_0 : 3'h0;
  assign v_10084_0 = v_601_0 ? v_3938_0 : 3'h0;
  assign v_10085_0 = v_10086_0 | v_10087_0;
  assign v_10086_0 = v_607_0 ? v_3952_0 : 3'h0;
  assign v_10087_0 = v_26_0 ? v_3938_0 : 3'h0;
  assign v_10088_0 = v_601_0 ? v_3931_0 : 3'h0;
  assign v_10089_0 = v_10090_0 | v_10091_0;
  assign v_10090_0 = v_607_0 ? v_3945_0 : 3'h0;
  assign v_10091_0 = v_26_0 ? v_3931_0 : 3'h0;
  assign v_10092_0 = v_601_0 ? v_3924_0 : 3'h0;
  assign v_10093_0 = v_10094_0 | v_10095_0;
  assign v_10094_0 = v_607_0 ? v_3938_0 : 3'h0;
  assign v_10095_0 = v_26_0 ? v_3924_0 : 3'h0;
  assign v_10096_0 = v_601_0 ? v_3917_0 : 3'h0;
  assign v_10097_0 = v_10098_0 | v_10099_0;
  assign v_10098_0 = v_607_0 ? v_3931_0 : 3'h0;
  assign v_10099_0 = v_26_0 ? v_3917_0 : 3'h0;
  assign v_10100_0 = v_601_0 ? v_3910_0 : 3'h0;
  assign v_10101_0 = v_10102_0 | v_10103_0;
  assign v_10102_0 = v_607_0 ? v_3924_0 : 3'h0;
  assign v_10103_0 = v_26_0 ? v_3910_0 : 3'h0;
  assign v_10104_0 = v_601_0 ? v_3903_0 : 3'h0;
  assign v_10105_0 = v_10106_0 | v_10107_0;
  assign v_10106_0 = v_607_0 ? v_3917_0 : 3'h0;
  assign v_10107_0 = v_26_0 ? v_3903_0 : 3'h0;
  assign v_10108_0 = v_601_0 ? v_3896_0 : 3'h0;
  assign v_10109_0 = v_10110_0 | v_10111_0;
  assign v_10110_0 = v_607_0 ? v_3910_0 : 3'h0;
  assign v_10111_0 = v_26_0 ? v_3896_0 : 3'h0;
  assign v_10112_0 = v_601_0 ? v_3889_0 : 3'h0;
  assign v_10113_0 = v_10114_0 | v_10115_0;
  assign v_10114_0 = v_607_0 ? v_3903_0 : 3'h0;
  assign v_10115_0 = v_26_0 ? v_3889_0 : 3'h0;
  assign v_10116_0 = v_601_0 ? v_3882_0 : 3'h0;
  assign v_10117_0 = v_10118_0 | v_10119_0;
  assign v_10118_0 = v_607_0 ? v_3896_0 : 3'h0;
  assign v_10119_0 = v_26_0 ? v_3882_0 : 3'h0;
  assign v_10120_0 = v_601_0 ? v_3875_0 : 3'h0;
  assign v_10121_0 = v_10122_0 | v_10123_0;
  assign v_10122_0 = v_607_0 ? v_3889_0 : 3'h0;
  assign v_10123_0 = v_26_0 ? v_3875_0 : 3'h0;
  assign v_10124_0 = v_601_0 ? v_3868_0 : 3'h0;
  assign v_10125_0 = v_10126_0 | v_10127_0;
  assign v_10126_0 = v_607_0 ? v_3882_0 : 3'h0;
  assign v_10127_0 = v_26_0 ? v_3868_0 : 3'h0;
  assign v_10128_0 = v_601_0 ? v_3861_0 : 3'h0;
  assign v_10129_0 = v_10130_0 | v_10131_0;
  assign v_10130_0 = v_607_0 ? v_3875_0 : 3'h0;
  assign v_10131_0 = v_26_0 ? v_3861_0 : 3'h0;
  assign v_10132_0 = v_601_0 ? v_3854_0 : 3'h0;
  assign v_10133_0 = v_10134_0 | v_10135_0;
  assign v_10134_0 = v_607_0 ? v_3868_0 : 3'h0;
  assign v_10135_0 = v_26_0 ? v_3854_0 : 3'h0;
  assign v_10136_0 = v_601_0 ? v_3847_0 : 3'h0;
  assign v_10137_0 = v_10138_0 | v_10139_0;
  assign v_10138_0 = v_607_0 ? v_3861_0 : 3'h0;
  assign v_10139_0 = v_26_0 ? v_3847_0 : 3'h0;
  assign v_10140_0 = v_601_0 ? v_3840_0 : 3'h0;
  assign v_10141_0 = v_10142_0 | v_10143_0;
  assign v_10142_0 = v_607_0 ? v_3854_0 : 3'h0;
  assign v_10143_0 = v_26_0 ? v_3840_0 : 3'h0;
  assign v_10144_0 = v_601_0 ? v_3833_0 : 3'h0;
  assign v_10145_0 = v_10146_0 | v_10147_0;
  assign v_10146_0 = v_607_0 ? v_3847_0 : 3'h0;
  assign v_10147_0 = v_26_0 ? v_3833_0 : 3'h0;
  assign v_10148_0 = v_601_0 ? v_3826_0 : 3'h0;
  assign v_10149_0 = v_10150_0 | v_10151_0;
  assign v_10150_0 = v_607_0 ? v_3840_0 : 3'h0;
  assign v_10151_0 = v_26_0 ? v_3826_0 : 3'h0;
  assign v_10152_0 = v_601_0 ? v_3819_0 : 3'h0;
  assign v_10153_0 = v_10154_0 | v_10155_0;
  assign v_10154_0 = v_607_0 ? v_3833_0 : 3'h0;
  assign v_10155_0 = v_26_0 ? v_3819_0 : 3'h0;
  assign v_10156_0 = v_601_0 ? v_3812_0 : 3'h0;
  assign v_10157_0 = v_10158_0 | v_10159_0;
  assign v_10158_0 = v_607_0 ? v_3826_0 : 3'h0;
  assign v_10159_0 = v_26_0 ? v_3812_0 : 3'h0;
  assign v_10160_0 = v_601_0 ? v_3805_0 : 3'h0;
  assign v_10161_0 = v_10162_0 | v_10163_0;
  assign v_10162_0 = v_607_0 ? v_3819_0 : 3'h0;
  assign v_10163_0 = v_26_0 ? v_3805_0 : 3'h0;
  assign v_10164_0 = v_601_0 ? v_3798_0 : 3'h0;
  assign v_10165_0 = v_10166_0 | v_10167_0;
  assign v_10166_0 = v_607_0 ? v_3812_0 : 3'h0;
  assign v_10167_0 = v_26_0 ? v_3798_0 : 3'h0;
  assign v_10168_0 = v_601_0 ? v_3791_0 : 3'h0;
  assign v_10169_0 = v_10170_0 | v_10171_0;
  assign v_10170_0 = v_607_0 ? v_3805_0 : 3'h0;
  assign v_10171_0 = v_26_0 ? v_3791_0 : 3'h0;
  assign v_10172_0 = v_601_0 ? v_3784_0 : 3'h0;
  assign v_10173_0 = v_10174_0 | v_10175_0;
  assign v_10174_0 = v_607_0 ? v_3798_0 : 3'h0;
  assign v_10175_0 = v_26_0 ? v_3784_0 : 3'h0;
  assign v_10176_0 = v_601_0 ? v_3777_0 : 3'h0;
  assign v_10177_0 = v_10178_0 | v_10179_0;
  assign v_10178_0 = v_607_0 ? v_3791_0 : 3'h0;
  assign v_10179_0 = v_26_0 ? v_3777_0 : 3'h0;
  assign v_10180_0 = v_601_0 ? v_3770_0 : 3'h0;
  assign v_10181_0 = v_10182_0 | v_10183_0;
  assign v_10182_0 = v_607_0 ? v_3784_0 : 3'h0;
  assign v_10183_0 = v_26_0 ? v_3770_0 : 3'h0;
  assign v_10184_0 = v_601_0 ? v_3763_0 : 3'h0;
  assign v_10185_0 = v_10186_0 | v_10187_0;
  assign v_10186_0 = v_607_0 ? v_3777_0 : 3'h0;
  assign v_10187_0 = v_26_0 ? v_3763_0 : 3'h0;
  assign v_10188_0 = v_601_0 ? v_3756_0 : 3'h0;
  assign v_10189_0 = v_10190_0 | v_10191_0;
  assign v_10190_0 = v_607_0 ? v_3770_0 : 3'h0;
  assign v_10191_0 = v_26_0 ? v_3756_0 : 3'h0;
  assign v_10192_0 = v_601_0 ? v_3749_0 : 3'h0;
  assign v_10193_0 = v_10194_0 | v_10195_0;
  assign v_10194_0 = v_607_0 ? v_3763_0 : 3'h0;
  assign v_10195_0 = v_26_0 ? v_3749_0 : 3'h0;
  assign v_10196_0 = v_601_0 ? v_3742_0 : 3'h0;
  assign v_10197_0 = v_10198_0 | v_10199_0;
  assign v_10198_0 = v_607_0 ? v_3756_0 : 3'h0;
  assign v_10199_0 = v_26_0 ? v_3742_0 : 3'h0;
  assign v_10200_0 = v_601_0 ? v_3735_0 : 3'h0;
  assign v_10201_0 = v_10202_0 | v_10203_0;
  assign v_10202_0 = v_607_0 ? v_3749_0 : 3'h0;
  assign v_10203_0 = v_26_0 ? v_3735_0 : 3'h0;
  assign v_10204_0 = v_601_0 ? v_3728_0 : 3'h0;
  assign v_10205_0 = v_10206_0 | v_10207_0;
  assign v_10206_0 = v_607_0 ? v_3742_0 : 3'h0;
  assign v_10207_0 = v_26_0 ? v_3728_0 : 3'h0;
  assign v_10208_0 = v_601_0 ? v_3721_0 : 3'h0;
  assign v_10209_0 = v_10210_0 | v_10211_0;
  assign v_10210_0 = v_607_0 ? v_3735_0 : 3'h0;
  assign v_10211_0 = v_26_0 ? v_3721_0 : 3'h0;
  assign v_10212_0 = v_601_0 ? v_3714_0 : 3'h0;
  assign v_10213_0 = v_10214_0 | v_10215_0;
  assign v_10214_0 = v_607_0 ? v_3728_0 : 3'h0;
  assign v_10215_0 = v_26_0 ? v_3714_0 : 3'h0;
  assign v_10216_0 = v_601_0 ? v_3707_0 : 3'h0;
  assign v_10217_0 = v_10218_0 | v_10219_0;
  assign v_10218_0 = v_607_0 ? v_3721_0 : 3'h0;
  assign v_10219_0 = v_26_0 ? v_3707_0 : 3'h0;
  assign v_10220_0 = v_601_0 ? v_3700_0 : 3'h0;
  assign v_10221_0 = v_10222_0 | v_10223_0;
  assign v_10222_0 = v_607_0 ? v_3714_0 : 3'h0;
  assign v_10223_0 = v_26_0 ? v_3700_0 : 3'h0;
  assign v_10224_0 = v_601_0 ? v_3693_0 : 3'h0;
  assign v_10225_0 = v_10226_0 | v_10227_0;
  assign v_10226_0 = v_607_0 ? v_3707_0 : 3'h0;
  assign v_10227_0 = v_26_0 ? v_3693_0 : 3'h0;
  assign v_10228_0 = v_601_0 ? v_3686_0 : 3'h0;
  assign v_10229_0 = v_10230_0 | v_10231_0;
  assign v_10230_0 = v_607_0 ? v_3700_0 : 3'h0;
  assign v_10231_0 = v_26_0 ? v_3686_0 : 3'h0;
  assign v_10232_0 = v_601_0 ? v_3679_0 : 3'h0;
  assign v_10233_0 = v_10234_0 | v_10235_0;
  assign v_10234_0 = v_607_0 ? v_3693_0 : 3'h0;
  assign v_10235_0 = v_26_0 ? v_3679_0 : 3'h0;
  assign v_10236_0 = v_601_0 ? v_3672_0 : 3'h0;
  assign v_10237_0 = v_10238_0 | v_10239_0;
  assign v_10238_0 = v_607_0 ? v_3686_0 : 3'h0;
  assign v_10239_0 = v_26_0 ? v_3672_0 : 3'h0;
  assign v_10240_0 = v_601_0 ? v_3665_0 : 3'h0;
  assign v_10241_0 = v_10242_0 | v_10243_0;
  assign v_10242_0 = v_607_0 ? v_3679_0 : 3'h0;
  assign v_10243_0 = v_26_0 ? v_3665_0 : 3'h0;
  assign v_10244_0 = v_601_0 ? v_3658_0 : 3'h0;
  assign v_10245_0 = v_10246_0 | v_10247_0;
  assign v_10246_0 = v_607_0 ? v_3672_0 : 3'h0;
  assign v_10247_0 = v_26_0 ? v_3658_0 : 3'h0;
  assign v_10248_0 = v_601_0 ? v_3651_0 : 3'h0;
  assign v_10249_0 = v_10250_0 | v_10251_0;
  assign v_10250_0 = v_607_0 ? v_3665_0 : 3'h0;
  assign v_10251_0 = v_26_0 ? v_3651_0 : 3'h0;
  assign v_10252_0 = v_601_0 ? v_3644_0 : 3'h0;
  assign v_10253_0 = v_10254_0 | v_10255_0;
  assign v_10254_0 = v_607_0 ? v_3658_0 : 3'h0;
  assign v_10255_0 = v_26_0 ? v_3644_0 : 3'h0;
  assign v_10256_0 = v_601_0 ? v_3637_0 : 3'h0;
  assign v_10257_0 = v_10258_0 | v_10259_0;
  assign v_10258_0 = v_607_0 ? v_3651_0 : 3'h0;
  assign v_10259_0 = v_26_0 ? v_3637_0 : 3'h0;
  assign v_10260_0 = v_601_0 ? v_3630_0 : 3'h0;
  assign v_10261_0 = v_10262_0 | v_10263_0;
  assign v_10262_0 = v_607_0 ? v_3644_0 : 3'h0;
  assign v_10263_0 = v_26_0 ? v_3630_0 : 3'h0;
  assign v_10264_0 = v_601_0 ? v_3623_0 : 3'h0;
  assign v_10265_0 = v_10266_0 | v_10267_0;
  assign v_10266_0 = v_607_0 ? v_3637_0 : 3'h0;
  assign v_10267_0 = v_26_0 ? v_3623_0 : 3'h0;
  assign v_10268_0 = v_601_0 ? v_3616_0 : 3'h0;
  assign v_10269_0 = v_10270_0 | v_10271_0;
  assign v_10270_0 = v_607_0 ? v_3630_0 : 3'h0;
  assign v_10271_0 = v_26_0 ? v_3616_0 : 3'h0;
  assign v_10272_0 = v_601_0 ? v_3609_0 : 3'h0;
  assign v_10273_0 = v_10274_0 | v_10275_0;
  assign v_10274_0 = v_607_0 ? v_3623_0 : 3'h0;
  assign v_10275_0 = v_26_0 ? v_3609_0 : 3'h0;
  assign v_10276_0 = v_601_0 ? v_3602_0 : 3'h0;
  assign v_10277_0 = v_10278_0 | v_10279_0;
  assign v_10278_0 = v_607_0 ? v_3616_0 : 3'h0;
  assign v_10279_0 = v_26_0 ? v_3602_0 : 3'h0;
  assign v_10280_0 = v_601_0 ? v_3595_0 : 3'h0;
  assign v_10281_0 = v_10282_0 | v_10283_0;
  assign v_10282_0 = v_607_0 ? v_3609_0 : 3'h0;
  assign v_10283_0 = v_26_0 ? v_3595_0 : 3'h0;
  assign v_10284_0 = v_601_0 ? v_3588_0 : 3'h0;
  assign v_10285_0 = v_10286_0 | v_10287_0;
  assign v_10286_0 = v_607_0 ? v_3602_0 : 3'h0;
  assign v_10287_0 = v_26_0 ? v_3588_0 : 3'h0;
  assign v_10288_0 = v_601_0 ? v_3581_0 : 3'h0;
  assign v_10289_0 = v_10290_0 | v_10291_0;
  assign v_10290_0 = v_607_0 ? v_3595_0 : 3'h0;
  assign v_10291_0 = v_26_0 ? v_3581_0 : 3'h0;
  assign v_10292_0 = v_601_0 ? v_3574_0 : 3'h0;
  assign v_10293_0 = v_10294_0 | v_10295_0;
  assign v_10294_0 = v_607_0 ? v_3588_0 : 3'h0;
  assign v_10295_0 = v_26_0 ? v_3574_0 : 3'h0;
  assign v_10296_0 = v_601_0 ? v_3567_0 : 3'h0;
  assign v_10297_0 = v_10298_0 | v_10299_0;
  assign v_10298_0 = v_607_0 ? v_3581_0 : 3'h0;
  assign v_10299_0 = v_26_0 ? v_3567_0 : 3'h0;
  assign v_10300_0 = v_601_0 ? v_3560_0 : 3'h0;
  assign v_10301_0 = v_10302_0 | v_10303_0;
  assign v_10302_0 = v_607_0 ? v_3574_0 : 3'h0;
  assign v_10303_0 = v_26_0 ? v_3560_0 : 3'h0;
  assign v_10304_0 = v_601_0 ? v_3553_0 : 3'h0;
  assign v_10305_0 = v_10306_0 | v_10307_0;
  assign v_10306_0 = v_607_0 ? v_3567_0 : 3'h0;
  assign v_10307_0 = v_26_0 ? v_3553_0 : 3'h0;
  assign v_10308_0 = v_601_0 ? v_3546_0 : 3'h0;
  assign v_10309_0 = v_10310_0 | v_10311_0;
  assign v_10310_0 = v_607_0 ? v_3560_0 : 3'h0;
  assign v_10311_0 = v_26_0 ? v_3546_0 : 3'h0;
  assign v_10312_0 = v_601_0 ? v_3539_0 : 3'h0;
  assign v_10313_0 = v_10314_0 | v_10315_0;
  assign v_10314_0 = v_607_0 ? v_3553_0 : 3'h0;
  assign v_10315_0 = v_26_0 ? v_3539_0 : 3'h0;
  assign v_10316_0 = v_601_0 ? v_3532_0 : 3'h0;
  assign v_10317_0 = v_10318_0 | v_10319_0;
  assign v_10318_0 = v_607_0 ? v_3546_0 : 3'h0;
  assign v_10319_0 = v_26_0 ? v_3532_0 : 3'h0;
  assign v_10320_0 = v_601_0 ? v_3525_0 : 3'h0;
  assign v_10321_0 = v_10322_0 | v_10323_0;
  assign v_10322_0 = v_607_0 ? v_3539_0 : 3'h0;
  assign v_10323_0 = v_26_0 ? v_3525_0 : 3'h0;
  assign v_10324_0 = v_601_0 ? v_3518_0 : 3'h0;
  assign v_10325_0 = v_10326_0 | v_10327_0;
  assign v_10326_0 = v_607_0 ? v_3532_0 : 3'h0;
  assign v_10327_0 = v_26_0 ? v_3518_0 : 3'h0;
  assign v_10328_0 = v_601_0 ? v_3511_0 : 3'h0;
  assign v_10329_0 = v_10330_0 | v_10331_0;
  assign v_10330_0 = v_607_0 ? v_3525_0 : 3'h0;
  assign v_10331_0 = v_26_0 ? v_3511_0 : 3'h0;
  assign v_10332_0 = v_601_0 ? v_3504_0 : 3'h0;
  assign v_10333_0 = v_10334_0 | v_10335_0;
  assign v_10334_0 = v_607_0 ? v_3518_0 : 3'h0;
  assign v_10335_0 = v_26_0 ? v_3504_0 : 3'h0;
  assign v_10336_0 = v_601_0 ? v_3497_0 : 3'h0;
  assign v_10337_0 = v_10338_0 | v_10339_0;
  assign v_10338_0 = v_607_0 ? v_3511_0 : 3'h0;
  assign v_10339_0 = v_26_0 ? v_3497_0 : 3'h0;
  assign v_10340_0 = v_601_0 ? v_3490_0 : 3'h0;
  assign v_10341_0 = v_10342_0 | v_10343_0;
  assign v_10342_0 = v_607_0 ? v_3504_0 : 3'h0;
  assign v_10343_0 = v_26_0 ? v_3490_0 : 3'h0;
  assign v_10344_0 = v_601_0 ? v_3483_0 : 3'h0;
  assign v_10345_0 = v_10346_0 | v_10347_0;
  assign v_10346_0 = v_607_0 ? v_3497_0 : 3'h0;
  assign v_10347_0 = v_26_0 ? v_3483_0 : 3'h0;
  assign v_10348_0 = v_601_0 ? v_3476_0 : 3'h0;
  assign v_10349_0 = v_10350_0 | v_10351_0;
  assign v_10350_0 = v_607_0 ? v_3490_0 : 3'h0;
  assign v_10351_0 = v_26_0 ? v_3476_0 : 3'h0;
  assign v_10352_0 = v_601_0 ? v_3469_0 : 3'h0;
  assign v_10353_0 = v_10354_0 | v_10355_0;
  assign v_10354_0 = v_607_0 ? v_3483_0 : 3'h0;
  assign v_10355_0 = v_26_0 ? v_3469_0 : 3'h0;
  assign v_10356_0 = v_601_0 ? v_3462_0 : 3'h0;
  assign v_10357_0 = v_10358_0 | v_10359_0;
  assign v_10358_0 = v_607_0 ? v_3476_0 : 3'h0;
  assign v_10359_0 = v_26_0 ? v_3462_0 : 3'h0;
  assign v_10360_0 = v_601_0 ? v_3455_0 : 3'h0;
  assign v_10361_0 = v_10362_0 | v_10363_0;
  assign v_10362_0 = v_607_0 ? v_3469_0 : 3'h0;
  assign v_10363_0 = v_26_0 ? v_3455_0 : 3'h0;
  assign v_10364_0 = v_601_0 ? v_3448_0 : 3'h0;
  assign v_10365_0 = v_10366_0 | v_10367_0;
  assign v_10366_0 = v_607_0 ? v_3462_0 : 3'h0;
  assign v_10367_0 = v_26_0 ? v_3448_0 : 3'h0;
  assign v_10368_0 = v_601_0 ? v_3441_0 : 3'h0;
  assign v_10369_0 = v_10370_0 | v_10371_0;
  assign v_10370_0 = v_607_0 ? v_3455_0 : 3'h0;
  assign v_10371_0 = v_26_0 ? v_3441_0 : 3'h0;
  assign v_10372_0 = v_601_0 ? v_3434_0 : 3'h0;
  assign v_10373_0 = v_10374_0 | v_10375_0;
  assign v_10374_0 = v_607_0 ? v_3448_0 : 3'h0;
  assign v_10375_0 = v_26_0 ? v_3434_0 : 3'h0;
  assign v_10376_0 = v_601_0 ? v_3427_0 : 3'h0;
  assign v_10377_0 = v_10378_0 | v_10379_0;
  assign v_10378_0 = v_607_0 ? v_3441_0 : 3'h0;
  assign v_10379_0 = v_26_0 ? v_3427_0 : 3'h0;
  assign v_10380_0 = v_601_0 ? v_3420_0 : 3'h0;
  assign v_10381_0 = v_10382_0 | v_10383_0;
  assign v_10382_0 = v_607_0 ? v_3434_0 : 3'h0;
  assign v_10383_0 = v_26_0 ? v_3420_0 : 3'h0;
  assign v_10384_0 = v_601_0 ? v_3413_0 : 3'h0;
  assign v_10385_0 = v_10386_0 | v_10387_0;
  assign v_10386_0 = v_607_0 ? v_3427_0 : 3'h0;
  assign v_10387_0 = v_26_0 ? v_3413_0 : 3'h0;
  assign v_10388_0 = v_601_0 ? v_3406_0 : 3'h0;
  assign v_10389_0 = v_10390_0 | v_10391_0;
  assign v_10390_0 = v_607_0 ? v_3420_0 : 3'h0;
  assign v_10391_0 = v_26_0 ? v_3406_0 : 3'h0;
  assign v_10392_0 = v_601_0 ? v_3399_0 : 3'h0;
  assign v_10393_0 = v_10394_0 | v_10395_0;
  assign v_10394_0 = v_607_0 ? v_3413_0 : 3'h0;
  assign v_10395_0 = v_26_0 ? v_3399_0 : 3'h0;
  assign v_10396_0 = v_601_0 ? v_3392_0 : 3'h0;
  assign v_10397_0 = v_10398_0 | v_10399_0;
  assign v_10398_0 = v_607_0 ? v_3406_0 : 3'h0;
  assign v_10399_0 = v_26_0 ? v_3392_0 : 3'h0;
  assign v_10400_0 = v_601_0 ? v_3385_0 : 3'h0;
  assign v_10401_0 = v_10402_0 | v_10403_0;
  assign v_10402_0 = v_607_0 ? v_3399_0 : 3'h0;
  assign v_10403_0 = v_26_0 ? v_3385_0 : 3'h0;
  assign v_10404_0 = v_601_0 ? v_3378_0 : 3'h0;
  assign v_10405_0 = v_10406_0 | v_10407_0;
  assign v_10406_0 = v_607_0 ? v_3392_0 : 3'h0;
  assign v_10407_0 = v_26_0 ? v_3378_0 : 3'h0;
  assign v_10408_0 = v_601_0 ? v_3371_0 : 3'h0;
  assign v_10409_0 = v_10410_0 | v_10411_0;
  assign v_10410_0 = v_607_0 ? v_3385_0 : 3'h0;
  assign v_10411_0 = v_26_0 ? v_3371_0 : 3'h0;
  assign v_10412_0 = v_601_0 ? v_3364_0 : 3'h0;
  assign v_10413_0 = v_10414_0 | v_10415_0;
  assign v_10414_0 = v_607_0 ? v_3378_0 : 3'h0;
  assign v_10415_0 = v_26_0 ? v_3364_0 : 3'h0;
  assign v_10416_0 = v_601_0 ? v_3357_0 : 3'h0;
  assign v_10417_0 = v_10418_0 | v_10419_0;
  assign v_10418_0 = v_607_0 ? v_3371_0 : 3'h0;
  assign v_10419_0 = v_26_0 ? v_3357_0 : 3'h0;
  assign v_10420_0 = v_601_0 ? v_3350_0 : 3'h0;
  assign v_10421_0 = v_10422_0 | v_10423_0;
  assign v_10422_0 = v_607_0 ? v_3364_0 : 3'h0;
  assign v_10423_0 = v_26_0 ? v_3350_0 : 3'h0;
  assign v_10424_0 = v_601_0 ? v_3343_0 : 3'h0;
  assign v_10425_0 = v_10426_0 | v_10427_0;
  assign v_10426_0 = v_607_0 ? v_3357_0 : 3'h0;
  assign v_10427_0 = v_26_0 ? v_3343_0 : 3'h0;
  assign v_10428_0 = v_601_0 ? v_3336_0 : 3'h0;
  assign v_10429_0 = v_10430_0 | v_10431_0;
  assign v_10430_0 = v_607_0 ? v_3350_0 : 3'h0;
  assign v_10431_0 = v_26_0 ? v_3336_0 : 3'h0;
  assign v_10432_0 = v_601_0 ? v_3329_0 : 3'h0;
  assign v_10433_0 = v_10434_0 | v_10435_0;
  assign v_10434_0 = v_607_0 ? v_3343_0 : 3'h0;
  assign v_10435_0 = v_26_0 ? v_3329_0 : 3'h0;
  assign v_10436_0 = v_601_0 ? v_3322_0 : 3'h0;
  assign v_10437_0 = v_10438_0 | v_10439_0;
  assign v_10438_0 = v_607_0 ? v_3336_0 : 3'h0;
  assign v_10439_0 = v_26_0 ? v_3322_0 : 3'h0;
  assign v_10440_0 = v_601_0 ? v_3315_0 : 3'h0;
  assign v_10441_0 = v_10442_0 | v_10443_0;
  assign v_10442_0 = v_607_0 ? v_3329_0 : 3'h0;
  assign v_10443_0 = v_26_0 ? v_3315_0 : 3'h0;
  assign v_10444_0 = v_601_0 ? v_3308_0 : 3'h0;
  assign v_10445_0 = v_10446_0 | v_10447_0;
  assign v_10446_0 = v_607_0 ? v_3322_0 : 3'h0;
  assign v_10447_0 = v_26_0 ? v_3308_0 : 3'h0;
  assign v_10448_0 = v_601_0 ? v_3301_0 : 3'h0;
  assign v_10449_0 = v_10450_0 | v_10451_0;
  assign v_10450_0 = v_607_0 ? v_3315_0 : 3'h0;
  assign v_10451_0 = v_26_0 ? v_3301_0 : 3'h0;
  assign v_10452_0 = v_601_0 ? v_3294_0 : 3'h0;
  assign v_10453_0 = v_10454_0 | v_10455_0;
  assign v_10454_0 = v_607_0 ? v_3308_0 : 3'h0;
  assign v_10455_0 = v_26_0 ? v_3294_0 : 3'h0;
  assign v_10456_0 = v_601_0 ? v_3287_0 : 3'h0;
  assign v_10457_0 = v_10458_0 | v_10459_0;
  assign v_10458_0 = v_607_0 ? v_3301_0 : 3'h0;
  assign v_10459_0 = v_26_0 ? v_3287_0 : 3'h0;
  assign v_10460_0 = v_601_0 ? v_3280_0 : 3'h0;
  assign v_10461_0 = v_10462_0 | v_10463_0;
  assign v_10462_0 = v_607_0 ? v_3294_0 : 3'h0;
  assign v_10463_0 = v_26_0 ? v_3280_0 : 3'h0;
  assign v_10464_0 = v_601_0 ? v_3273_0 : 3'h0;
  assign v_10465_0 = v_10466_0 | v_10467_0;
  assign v_10466_0 = v_607_0 ? v_3287_0 : 3'h0;
  assign v_10467_0 = v_26_0 ? v_3273_0 : 3'h0;
  assign v_10468_0 = v_601_0 ? v_3266_0 : 3'h0;
  assign v_10469_0 = v_10470_0 | v_10471_0;
  assign v_10470_0 = v_607_0 ? v_3280_0 : 3'h0;
  assign v_10471_0 = v_26_0 ? v_3266_0 : 3'h0;
  assign v_10472_0 = v_601_0 ? v_3259_0 : 3'h0;
  assign v_10473_0 = v_10474_0 | v_10475_0;
  assign v_10474_0 = v_607_0 ? v_3273_0 : 3'h0;
  assign v_10475_0 = v_26_0 ? v_3259_0 : 3'h0;
  assign v_10476_0 = v_601_0 ? v_3252_0 : 3'h0;
  assign v_10477_0 = v_10478_0 | v_10479_0;
  assign v_10478_0 = v_607_0 ? v_3266_0 : 3'h0;
  assign v_10479_0 = v_26_0 ? v_3252_0 : 3'h0;
  assign v_10480_0 = v_601_0 ? v_3245_0 : 3'h0;
  assign v_10481_0 = v_10482_0 | v_10483_0;
  assign v_10482_0 = v_607_0 ? v_3259_0 : 3'h0;
  assign v_10483_0 = v_26_0 ? v_3245_0 : 3'h0;
  assign v_10484_0 = v_601_0 ? v_3238_0 : 3'h0;
  assign v_10485_0 = v_10486_0 | v_10487_0;
  assign v_10486_0 = v_607_0 ? v_3252_0 : 3'h0;
  assign v_10487_0 = v_26_0 ? v_3238_0 : 3'h0;
  assign v_10488_0 = v_601_0 ? v_3231_0 : 3'h0;
  assign v_10489_0 = v_10490_0 | v_10491_0;
  assign v_10490_0 = v_607_0 ? v_3245_0 : 3'h0;
  assign v_10491_0 = v_26_0 ? v_3231_0 : 3'h0;
  assign v_10492_0 = v_601_0 ? v_3224_0 : 3'h0;
  assign v_10493_0 = v_10494_0 | v_10495_0;
  assign v_10494_0 = v_607_0 ? v_3238_0 : 3'h0;
  assign v_10495_0 = v_26_0 ? v_3224_0 : 3'h0;
  assign v_10496_0 = v_601_0 ? v_3217_0 : 3'h0;
  assign v_10497_0 = v_10498_0 | v_10499_0;
  assign v_10498_0 = v_607_0 ? v_3231_0 : 3'h0;
  assign v_10499_0 = v_26_0 ? v_3217_0 : 3'h0;
  assign v_10500_0 = v_601_0 ? v_3210_0 : 3'h0;
  assign v_10501_0 = v_10502_0 | v_10503_0;
  assign v_10502_0 = v_607_0 ? v_3224_0 : 3'h0;
  assign v_10503_0 = v_26_0 ? v_3210_0 : 3'h0;
  assign v_10504_0 = v_601_0 ? v_3203_0 : 3'h0;
  assign v_10505_0 = v_10506_0 | v_10507_0;
  assign v_10506_0 = v_607_0 ? v_3217_0 : 3'h0;
  assign v_10507_0 = v_26_0 ? v_3203_0 : 3'h0;
  assign v_10508_0 = v_601_0 ? v_3196_0 : 3'h0;
  assign v_10509_0 = v_10510_0 | v_10511_0;
  assign v_10510_0 = v_607_0 ? v_3210_0 : 3'h0;
  assign v_10511_0 = v_26_0 ? v_3196_0 : 3'h0;
  assign v_10512_0 = v_601_0 ? v_3189_0 : 3'h0;
  assign v_10513_0 = v_10514_0 | v_10515_0;
  assign v_10514_0 = v_607_0 ? v_3203_0 : 3'h0;
  assign v_10515_0 = v_26_0 ? v_3189_0 : 3'h0;
  assign v_10516_0 = v_601_0 ? v_3182_0 : 3'h0;
  assign v_10517_0 = v_10518_0 | v_10519_0;
  assign v_10518_0 = v_607_0 ? v_3196_0 : 3'h0;
  assign v_10519_0 = v_26_0 ? v_3182_0 : 3'h0;
  assign v_10520_0 = v_601_0 ? v_3175_0 : 3'h0;
  assign v_10521_0 = v_10522_0 | v_10523_0;
  assign v_10522_0 = v_607_0 ? v_3189_0 : 3'h0;
  assign v_10523_0 = v_26_0 ? v_3175_0 : 3'h0;
  assign v_10524_0 = v_601_0 ? v_3168_0 : 3'h0;
  assign v_10525_0 = v_10526_0 | v_10527_0;
  assign v_10526_0 = v_607_0 ? v_3182_0 : 3'h0;
  assign v_10527_0 = v_26_0 ? v_3168_0 : 3'h0;
  assign v_10528_0 = v_601_0 ? v_3161_0 : 3'h0;
  assign v_10529_0 = v_10530_0 | v_10531_0;
  assign v_10530_0 = v_607_0 ? v_3175_0 : 3'h0;
  assign v_10531_0 = v_26_0 ? v_3161_0 : 3'h0;
  assign v_10532_0 = v_601_0 ? v_3154_0 : 3'h0;
  assign v_10533_0 = v_10534_0 | v_10535_0;
  assign v_10534_0 = v_607_0 ? v_3168_0 : 3'h0;
  assign v_10535_0 = v_26_0 ? v_3154_0 : 3'h0;
  assign v_10536_0 = v_601_0 ? v_3147_0 : 3'h0;
  assign v_10537_0 = v_10538_0 | v_10539_0;
  assign v_10538_0 = v_607_0 ? v_3161_0 : 3'h0;
  assign v_10539_0 = v_26_0 ? v_3147_0 : 3'h0;
  assign v_10540_0 = v_601_0 ? v_3140_0 : 3'h0;
  assign v_10541_0 = v_10542_0 | v_10543_0;
  assign v_10542_0 = v_607_0 ? v_3154_0 : 3'h0;
  assign v_10543_0 = v_26_0 ? v_3140_0 : 3'h0;
  assign v_10544_0 = v_601_0 ? v_3133_0 : 3'h0;
  assign v_10545_0 = v_10546_0 | v_10547_0;
  assign v_10546_0 = v_607_0 ? v_3147_0 : 3'h0;
  assign v_10547_0 = v_26_0 ? v_3133_0 : 3'h0;
  assign v_10548_0 = v_601_0 ? v_3126_0 : 3'h0;
  assign v_10549_0 = v_10550_0 | v_10551_0;
  assign v_10550_0 = v_607_0 ? v_3140_0 : 3'h0;
  assign v_10551_0 = v_26_0 ? v_3126_0 : 3'h0;
  assign v_10552_0 = v_601_0 ? v_3119_0 : 3'h0;
  assign v_10553_0 = v_10554_0 | v_10555_0;
  assign v_10554_0 = v_607_0 ? v_3133_0 : 3'h0;
  assign v_10555_0 = v_26_0 ? v_3119_0 : 3'h0;
  assign v_10556_0 = v_601_0 ? v_3112_0 : 3'h0;
  assign v_10557_0 = v_10558_0 | v_10559_0;
  assign v_10558_0 = v_607_0 ? v_3126_0 : 3'h0;
  assign v_10559_0 = v_26_0 ? v_3112_0 : 3'h0;
  assign v_10560_0 = v_601_0 ? v_3105_0 : 3'h0;
  assign v_10561_0 = v_10562_0 | v_10563_0;
  assign v_10562_0 = v_607_0 ? v_3119_0 : 3'h0;
  assign v_10563_0 = v_26_0 ? v_3105_0 : 3'h0;
  assign v_10564_0 = v_601_0 ? v_3098_0 : 3'h0;
  assign v_10565_0 = v_10566_0 | v_10567_0;
  assign v_10566_0 = v_607_0 ? v_3112_0 : 3'h0;
  assign v_10567_0 = v_26_0 ? v_3098_0 : 3'h0;
  assign v_10568_0 = v_601_0 ? v_3091_0 : 3'h0;
  assign v_10569_0 = v_10570_0 | v_10571_0;
  assign v_10570_0 = v_607_0 ? v_3105_0 : 3'h0;
  assign v_10571_0 = v_26_0 ? v_3091_0 : 3'h0;
  assign v_10572_0 = v_601_0 ? v_3084_0 : 3'h0;
  assign v_10573_0 = v_10574_0 | v_10575_0;
  assign v_10574_0 = v_607_0 ? v_3098_0 : 3'h0;
  assign v_10575_0 = v_26_0 ? v_3084_0 : 3'h0;
  assign v_10576_0 = v_601_0 ? v_3077_0 : 3'h0;
  assign v_10577_0 = v_10578_0 | v_10579_0;
  assign v_10578_0 = v_607_0 ? v_3091_0 : 3'h0;
  assign v_10579_0 = v_26_0 ? v_3077_0 : 3'h0;
  assign v_10580_0 = v_601_0 ? v_3070_0 : 3'h0;
  assign v_10581_0 = v_10582_0 | v_10583_0;
  assign v_10582_0 = v_607_0 ? v_3084_0 : 3'h0;
  assign v_10583_0 = v_26_0 ? v_3070_0 : 3'h0;
  assign v_10584_0 = v_601_0 ? v_3063_0 : 3'h0;
  assign v_10585_0 = v_10586_0 | v_10587_0;
  assign v_10586_0 = v_607_0 ? v_3077_0 : 3'h0;
  assign v_10587_0 = v_26_0 ? v_3063_0 : 3'h0;
  assign v_10588_0 = v_601_0 ? v_3056_0 : 3'h0;
  assign v_10589_0 = v_10590_0 | v_10591_0;
  assign v_10590_0 = v_607_0 ? v_3070_0 : 3'h0;
  assign v_10591_0 = v_26_0 ? v_3056_0 : 3'h0;
  assign v_10592_0 = v_601_0 ? v_3049_0 : 3'h0;
  assign v_10593_0 = v_10594_0 | v_10595_0;
  assign v_10594_0 = v_607_0 ? v_3063_0 : 3'h0;
  assign v_10595_0 = v_26_0 ? v_3049_0 : 3'h0;
  assign v_10596_0 = v_601_0 ? v_3042_0 : 3'h0;
  assign v_10597_0 = v_10598_0 | v_10599_0;
  assign v_10598_0 = v_607_0 ? v_3056_0 : 3'h0;
  assign v_10599_0 = v_26_0 ? v_3042_0 : 3'h0;
  assign v_10600_0 = v_601_0 ? v_3035_0 : 3'h0;
  assign v_10601_0 = v_10602_0 | v_10603_0;
  assign v_10602_0 = v_607_0 ? v_3049_0 : 3'h0;
  assign v_10603_0 = v_26_0 ? v_3035_0 : 3'h0;
  assign v_10604_0 = v_601_0 ? v_3028_0 : 3'h0;
  assign v_10605_0 = v_10606_0 | v_10607_0;
  assign v_10606_0 = v_607_0 ? v_3042_0 : 3'h0;
  assign v_10607_0 = v_26_0 ? v_3028_0 : 3'h0;
  assign v_10608_0 = v_601_0 ? v_3021_0 : 3'h0;
  assign v_10609_0 = v_10610_0 | v_10611_0;
  assign v_10610_0 = v_607_0 ? v_3035_0 : 3'h0;
  assign v_10611_0 = v_26_0 ? v_3021_0 : 3'h0;
  assign v_10612_0 = v_601_0 ? v_3014_0 : 3'h0;
  assign v_10613_0 = v_10614_0 | v_10615_0;
  assign v_10614_0 = v_607_0 ? v_3028_0 : 3'h0;
  assign v_10615_0 = v_26_0 ? v_3014_0 : 3'h0;
  assign v_10616_0 = v_601_0 ? v_3007_0 : 3'h0;
  assign v_10617_0 = v_10618_0 | v_10619_0;
  assign v_10618_0 = v_607_0 ? v_3021_0 : 3'h0;
  assign v_10619_0 = v_26_0 ? v_3007_0 : 3'h0;
  assign v_10620_0 = v_601_0 ? v_3000_0 : 3'h0;
  assign v_10621_0 = v_10622_0 | v_10623_0;
  assign v_10622_0 = v_607_0 ? v_3014_0 : 3'h0;
  assign v_10623_0 = v_26_0 ? v_3000_0 : 3'h0;
  assign v_10624_0 = v_601_0 ? v_2993_0 : 3'h0;
  assign v_10625_0 = v_10626_0 | v_10627_0;
  assign v_10626_0 = v_607_0 ? v_3007_0 : 3'h0;
  assign v_10627_0 = v_26_0 ? v_2993_0 : 3'h0;
  assign v_10628_0 = v_601_0 ? v_2986_0 : 3'h0;
  assign v_10629_0 = v_10630_0 | v_10631_0;
  assign v_10630_0 = v_607_0 ? v_3000_0 : 3'h0;
  assign v_10631_0 = v_26_0 ? v_2986_0 : 3'h0;
  assign v_10632_0 = v_601_0 ? v_2979_0 : 3'h0;
  assign v_10633_0 = v_10634_0 | v_10635_0;
  assign v_10634_0 = v_607_0 ? v_2993_0 : 3'h0;
  assign v_10635_0 = v_26_0 ? v_2979_0 : 3'h0;
  assign v_10636_0 = v_601_0 ? v_2972_0 : 3'h0;
  assign v_10637_0 = v_10638_0 | v_10639_0;
  assign v_10638_0 = v_607_0 ? v_2986_0 : 3'h0;
  assign v_10639_0 = v_26_0 ? v_2972_0 : 3'h0;
  assign v_10640_0 = v_601_0 ? v_2965_0 : 3'h0;
  assign v_10641_0 = v_10642_0 | v_10643_0;
  assign v_10642_0 = v_607_0 ? v_2979_0 : 3'h0;
  assign v_10643_0 = v_26_0 ? v_2965_0 : 3'h0;
  assign v_10644_0 = v_601_0 ? v_2958_0 : 3'h0;
  assign v_10645_0 = v_10646_0 | v_10647_0;
  assign v_10646_0 = v_607_0 ? v_2972_0 : 3'h0;
  assign v_10647_0 = v_26_0 ? v_2958_0 : 3'h0;
  assign v_10648_0 = v_601_0 ? v_2951_0 : 3'h0;
  assign v_10649_0 = v_10650_0 | v_10651_0;
  assign v_10650_0 = v_607_0 ? v_2965_0 : 3'h0;
  assign v_10651_0 = v_26_0 ? v_2951_0 : 3'h0;
  assign v_10652_0 = v_601_0 ? v_2944_0 : 3'h0;
  assign v_10653_0 = v_10654_0 | v_10655_0;
  assign v_10654_0 = v_607_0 ? v_2958_0 : 3'h0;
  assign v_10655_0 = v_26_0 ? v_2944_0 : 3'h0;
  assign v_10656_0 = v_601_0 ? v_2937_0 : 3'h0;
  assign v_10657_0 = v_10658_0 | v_10659_0;
  assign v_10658_0 = v_607_0 ? v_2951_0 : 3'h0;
  assign v_10659_0 = v_26_0 ? v_2937_0 : 3'h0;
  assign v_10660_0 = v_601_0 ? v_2930_0 : 3'h0;
  assign v_10661_0 = v_10662_0 | v_10663_0;
  assign v_10662_0 = v_607_0 ? v_2944_0 : 3'h0;
  assign v_10663_0 = v_26_0 ? v_2930_0 : 3'h0;
  assign v_10664_0 = v_601_0 ? v_2923_0 : 3'h0;
  assign v_10665_0 = v_10666_0 | v_10667_0;
  assign v_10666_0 = v_607_0 ? v_2937_0 : 3'h0;
  assign v_10667_0 = v_26_0 ? v_2923_0 : 3'h0;
  assign v_10668_0 = v_601_0 ? v_2916_0 : 3'h0;
  assign v_10669_0 = v_10670_0 | v_10671_0;
  assign v_10670_0 = v_607_0 ? v_2930_0 : 3'h0;
  assign v_10671_0 = v_26_0 ? v_2916_0 : 3'h0;
  assign v_10672_0 = v_601_0 ? v_2909_0 : 3'h0;
  assign v_10673_0 = v_10674_0 | v_10675_0;
  assign v_10674_0 = v_607_0 ? v_2923_0 : 3'h0;
  assign v_10675_0 = v_26_0 ? v_2909_0 : 3'h0;
  assign v_10676_0 = v_601_0 ? v_2902_0 : 3'h0;
  assign v_10677_0 = v_10678_0 | v_10679_0;
  assign v_10678_0 = v_607_0 ? v_2916_0 : 3'h0;
  assign v_10679_0 = v_26_0 ? v_2902_0 : 3'h0;
  assign v_10680_0 = v_601_0 ? v_2895_0 : 3'h0;
  assign v_10681_0 = v_10682_0 | v_10683_0;
  assign v_10682_0 = v_607_0 ? v_2909_0 : 3'h0;
  assign v_10683_0 = v_26_0 ? v_2895_0 : 3'h0;
  assign v_10684_0 = v_601_0 ? v_2888_0 : 3'h0;
  assign v_10685_0 = v_10686_0 | v_10687_0;
  assign v_10686_0 = v_607_0 ? v_2902_0 : 3'h0;
  assign v_10687_0 = v_26_0 ? v_2888_0 : 3'h0;
  assign v_10688_0 = v_601_0 ? v_2881_0 : 3'h0;
  assign v_10689_0 = v_10690_0 | v_10691_0;
  assign v_10690_0 = v_607_0 ? v_2895_0 : 3'h0;
  assign v_10691_0 = v_26_0 ? v_2881_0 : 3'h0;
  assign v_10692_0 = v_601_0 ? v_2874_0 : 3'h0;
  assign v_10693_0 = v_10694_0 | v_10695_0;
  assign v_10694_0 = v_607_0 ? v_2888_0 : 3'h0;
  assign v_10695_0 = v_26_0 ? v_2874_0 : 3'h0;
  assign v_10696_0 = v_601_0 ? v_2867_0 : 3'h0;
  assign v_10697_0 = v_10698_0 | v_10699_0;
  assign v_10698_0 = v_607_0 ? v_2881_0 : 3'h0;
  assign v_10699_0 = v_26_0 ? v_2867_0 : 3'h0;
  assign v_10700_0 = v_601_0 ? v_2860_0 : 3'h0;
  assign v_10701_0 = v_10702_0 | v_10703_0;
  assign v_10702_0 = v_607_0 ? v_2874_0 : 3'h0;
  assign v_10703_0 = v_26_0 ? v_2860_0 : 3'h0;
  assign v_10704_0 = v_601_0 ? v_2853_0 : 3'h0;
  assign v_10705_0 = v_10706_0 | v_10707_0;
  assign v_10706_0 = v_607_0 ? v_2867_0 : 3'h0;
  assign v_10707_0 = v_26_0 ? v_2853_0 : 3'h0;
  assign v_10708_0 = v_601_0 ? v_2846_0 : 3'h0;
  assign v_10709_0 = v_10710_0 | v_10711_0;
  assign v_10710_0 = v_607_0 ? v_2860_0 : 3'h0;
  assign v_10711_0 = v_26_0 ? v_2846_0 : 3'h0;
  assign v_10712_0 = v_601_0 ? v_2839_0 : 3'h0;
  assign v_10713_0 = v_10714_0 | v_10715_0;
  assign v_10714_0 = v_607_0 ? v_2853_0 : 3'h0;
  assign v_10715_0 = v_26_0 ? v_2839_0 : 3'h0;
  assign v_10716_0 = v_601_0 ? v_2832_0 : 3'h0;
  assign v_10717_0 = v_10718_0 | v_10719_0;
  assign v_10718_0 = v_607_0 ? v_2846_0 : 3'h0;
  assign v_10719_0 = v_26_0 ? v_2832_0 : 3'h0;
  assign v_10720_0 = v_601_0 ? v_2825_0 : 3'h0;
  assign v_10721_0 = v_10722_0 | v_10723_0;
  assign v_10722_0 = v_607_0 ? v_2839_0 : 3'h0;
  assign v_10723_0 = v_26_0 ? v_2825_0 : 3'h0;
  assign v_10724_0 = v_601_0 ? v_2818_0 : 3'h0;
  assign v_10725_0 = v_10726_0 | v_10727_0;
  assign v_10726_0 = v_607_0 ? v_2832_0 : 3'h0;
  assign v_10727_0 = v_26_0 ? v_2818_0 : 3'h0;
  assign v_10728_0 = v_601_0 ? v_2811_0 : 3'h0;
  assign v_10729_0 = v_10730_0 | v_10731_0;
  assign v_10730_0 = v_607_0 ? v_2825_0 : 3'h0;
  assign v_10731_0 = v_26_0 ? v_2811_0 : 3'h0;
  assign v_10732_0 = v_601_0 ? v_2804_0 : 3'h0;
  assign v_10733_0 = v_10734_0 | v_10735_0;
  assign v_10734_0 = v_607_0 ? v_2818_0 : 3'h0;
  assign v_10735_0 = v_26_0 ? v_2804_0 : 3'h0;
  assign v_10736_0 = v_601_0 ? v_2797_0 : 3'h0;
  assign v_10737_0 = v_10738_0 | v_10739_0;
  assign v_10738_0 = v_607_0 ? v_2811_0 : 3'h0;
  assign v_10739_0 = v_26_0 ? v_2797_0 : 3'h0;
  assign v_10740_0 = v_601_0 ? v_2790_0 : 3'h0;
  assign v_10741_0 = v_10742_0 | v_10743_0;
  assign v_10742_0 = v_607_0 ? v_2804_0 : 3'h0;
  assign v_10743_0 = v_26_0 ? v_2790_0 : 3'h0;
  assign v_10744_0 = v_601_0 ? v_2783_0 : 3'h0;
  assign v_10745_0 = v_10746_0 | v_10747_0;
  assign v_10746_0 = v_607_0 ? v_2797_0 : 3'h0;
  assign v_10747_0 = v_26_0 ? v_2783_0 : 3'h0;
  assign v_10748_0 = v_601_0 ? v_2776_0 : 3'h0;
  assign v_10749_0 = v_10750_0 | v_10751_0;
  assign v_10750_0 = v_607_0 ? v_2790_0 : 3'h0;
  assign v_10751_0 = v_26_0 ? v_2776_0 : 3'h0;
  assign v_10752_0 = v_601_0 ? v_2769_0 : 3'h0;
  assign v_10753_0 = v_10754_0 | v_10755_0;
  assign v_10754_0 = v_607_0 ? v_2783_0 : 3'h0;
  assign v_10755_0 = v_26_0 ? v_2769_0 : 3'h0;
  assign v_10756_0 = v_601_0 ? v_2762_0 : 3'h0;
  assign v_10757_0 = v_10758_0 | v_10759_0;
  assign v_10758_0 = v_607_0 ? v_2776_0 : 3'h0;
  assign v_10759_0 = v_26_0 ? v_2762_0 : 3'h0;
  assign v_10760_0 = v_601_0 ? v_2755_0 : 3'h0;
  assign v_10761_0 = v_10762_0 | v_10763_0;
  assign v_10762_0 = v_607_0 ? v_2769_0 : 3'h0;
  assign v_10763_0 = v_26_0 ? v_2755_0 : 3'h0;
  assign v_10764_0 = v_601_0 ? v_2748_0 : 3'h0;
  assign v_10765_0 = v_10766_0 | v_10767_0;
  assign v_10766_0 = v_607_0 ? v_2762_0 : 3'h0;
  assign v_10767_0 = v_26_0 ? v_2748_0 : 3'h0;
  assign v_10768_0 = v_601_0 ? v_2741_0 : 3'h0;
  assign v_10769_0 = v_10770_0 | v_10771_0;
  assign v_10770_0 = v_607_0 ? v_2755_0 : 3'h0;
  assign v_10771_0 = v_26_0 ? v_2741_0 : 3'h0;
  assign v_10772_0 = v_601_0 ? v_2734_0 : 3'h0;
  assign v_10773_0 = v_10774_0 | v_10775_0;
  assign v_10774_0 = v_607_0 ? v_2748_0 : 3'h0;
  assign v_10775_0 = v_26_0 ? v_2734_0 : 3'h0;
  assign v_10776_0 = v_601_0 ? v_2727_0 : 3'h0;
  assign v_10777_0 = v_10778_0 | v_10779_0;
  assign v_10778_0 = v_607_0 ? v_2741_0 : 3'h0;
  assign v_10779_0 = v_26_0 ? v_2727_0 : 3'h0;
  assign v_10780_0 = v_601_0 ? v_2720_0 : 3'h0;
  assign v_10781_0 = v_10782_0 | v_10783_0;
  assign v_10782_0 = v_607_0 ? v_2734_0 : 3'h0;
  assign v_10783_0 = v_26_0 ? v_2720_0 : 3'h0;
  assign v_10784_0 = v_601_0 ? v_2713_0 : 3'h0;
  assign v_10785_0 = v_10786_0 | v_10787_0;
  assign v_10786_0 = v_607_0 ? v_2727_0 : 3'h0;
  assign v_10787_0 = v_26_0 ? v_2713_0 : 3'h0;
  assign v_10788_0 = v_601_0 ? v_2706_0 : 3'h0;
  assign v_10789_0 = v_10790_0 | v_10791_0;
  assign v_10790_0 = v_607_0 ? v_2720_0 : 3'h0;
  assign v_10791_0 = v_26_0 ? v_2706_0 : 3'h0;
  assign v_10792_0 = v_601_0 ? v_2699_0 : 3'h0;
  assign v_10793_0 = v_10794_0 | v_10795_0;
  assign v_10794_0 = v_607_0 ? v_2713_0 : 3'h0;
  assign v_10795_0 = v_26_0 ? v_2699_0 : 3'h0;
  assign v_10796_0 = v_601_0 ? v_2692_0 : 3'h0;
  assign v_10797_0 = v_10798_0 | v_10799_0;
  assign v_10798_0 = v_607_0 ? v_2706_0 : 3'h0;
  assign v_10799_0 = v_26_0 ? v_2692_0 : 3'h0;
  assign v_10800_0 = v_601_0 ? v_2685_0 : 3'h0;
  assign v_10801_0 = v_10802_0 | v_10803_0;
  assign v_10802_0 = v_607_0 ? v_2699_0 : 3'h0;
  assign v_10803_0 = v_26_0 ? v_2685_0 : 3'h0;
  assign v_10804_0 = v_601_0 ? v_2678_0 : 3'h0;
  assign v_10805_0 = v_10806_0 | v_10807_0;
  assign v_10806_0 = v_607_0 ? v_2692_0 : 3'h0;
  assign v_10807_0 = v_26_0 ? v_2678_0 : 3'h0;
  assign v_10808_0 = v_601_0 ? v_2671_0 : 3'h0;
  assign v_10809_0 = v_10810_0 | v_10811_0;
  assign v_10810_0 = v_607_0 ? v_2685_0 : 3'h0;
  assign v_10811_0 = v_26_0 ? v_2671_0 : 3'h0;
  assign v_10812_0 = v_601_0 ? v_2664_0 : 3'h0;
  assign v_10813_0 = v_10814_0 | v_10815_0;
  assign v_10814_0 = v_607_0 ? v_2678_0 : 3'h0;
  assign v_10815_0 = v_26_0 ? v_2664_0 : 3'h0;
  assign v_10816_0 = v_601_0 ? v_2657_0 : 3'h0;
  assign v_10817_0 = v_10818_0 | v_10819_0;
  assign v_10818_0 = v_607_0 ? v_2671_0 : 3'h0;
  assign v_10819_0 = v_26_0 ? v_2657_0 : 3'h0;
  assign v_10820_0 = v_601_0 ? v_2650_0 : 3'h0;
  assign v_10821_0 = v_10822_0 | v_10823_0;
  assign v_10822_0 = v_607_0 ? v_2664_0 : 3'h0;
  assign v_10823_0 = v_26_0 ? v_2650_0 : 3'h0;
  assign v_10824_0 = v_601_0 ? v_2643_0 : 3'h0;
  assign v_10825_0 = v_10826_0 | v_10827_0;
  assign v_10826_0 = v_607_0 ? v_2657_0 : 3'h0;
  assign v_10827_0 = v_26_0 ? v_2643_0 : 3'h0;
  assign v_10828_0 = v_601_0 ? v_2636_0 : 3'h0;
  assign v_10829_0 = v_10830_0 | v_10831_0;
  assign v_10830_0 = v_607_0 ? v_2650_0 : 3'h0;
  assign v_10831_0 = v_26_0 ? v_2636_0 : 3'h0;
  assign v_10832_0 = v_601_0 ? v_2629_0 : 3'h0;
  assign v_10833_0 = v_10834_0 | v_10835_0;
  assign v_10834_0 = v_607_0 ? v_2643_0 : 3'h0;
  assign v_10835_0 = v_26_0 ? v_2629_0 : 3'h0;
  assign v_10836_0 = v_601_0 ? v_2622_0 : 3'h0;
  assign v_10837_0 = v_10838_0 | v_10839_0;
  assign v_10838_0 = v_607_0 ? v_2636_0 : 3'h0;
  assign v_10839_0 = v_26_0 ? v_2622_0 : 3'h0;
  assign v_10840_0 = v_601_0 ? v_2615_0 : 3'h0;
  assign v_10841_0 = v_10842_0 | v_10843_0;
  assign v_10842_0 = v_607_0 ? v_2629_0 : 3'h0;
  assign v_10843_0 = v_26_0 ? v_2615_0 : 3'h0;
  assign v_10844_0 = v_601_0 ? v_2608_0 : 3'h0;
  assign v_10845_0 = v_10846_0 | v_10847_0;
  assign v_10846_0 = v_607_0 ? v_2622_0 : 3'h0;
  assign v_10847_0 = v_26_0 ? v_2608_0 : 3'h0;
  assign v_10848_0 = v_601_0 ? v_2601_0 : 3'h0;
  assign v_10849_0 = v_10850_0 | v_10851_0;
  assign v_10850_0 = v_607_0 ? v_2615_0 : 3'h0;
  assign v_10851_0 = v_26_0 ? v_2601_0 : 3'h0;
  assign v_10852_0 = v_601_0 ? v_2594_0 : 3'h0;
  assign v_10853_0 = v_10854_0 | v_10855_0;
  assign v_10854_0 = v_607_0 ? v_2608_0 : 3'h0;
  assign v_10855_0 = v_26_0 ? v_2594_0 : 3'h0;
  assign v_10856_0 = v_601_0 ? v_2587_0 : 3'h0;
  assign v_10857_0 = v_10858_0 | v_10859_0;
  assign v_10858_0 = v_607_0 ? v_2601_0 : 3'h0;
  assign v_10859_0 = v_26_0 ? v_2587_0 : 3'h0;
  assign v_10860_0 = v_601_0 ? v_2580_0 : 3'h0;
  assign v_10861_0 = v_10862_0 | v_10863_0;
  assign v_10862_0 = v_607_0 ? v_2594_0 : 3'h0;
  assign v_10863_0 = v_26_0 ? v_2580_0 : 3'h0;
  assign v_10864_0 = v_601_0 ? v_2573_0 : 3'h0;
  assign v_10865_0 = v_10866_0 | v_10867_0;
  assign v_10866_0 = v_607_0 ? v_2587_0 : 3'h0;
  assign v_10867_0 = v_26_0 ? v_2573_0 : 3'h0;
  assign v_10868_0 = v_601_0 ? v_2566_0 : 3'h0;
  assign v_10869_0 = v_10870_0 | v_10871_0;
  assign v_10870_0 = v_607_0 ? v_2580_0 : 3'h0;
  assign v_10871_0 = v_26_0 ? v_2566_0 : 3'h0;
  assign v_10872_0 = v_601_0 ? v_2559_0 : 3'h0;
  assign v_10873_0 = v_10874_0 | v_10875_0;
  assign v_10874_0 = v_607_0 ? v_2573_0 : 3'h0;
  assign v_10875_0 = v_26_0 ? v_2559_0 : 3'h0;
  assign v_10876_0 = v_601_0 ? v_2552_0 : 3'h0;
  assign v_10877_0 = v_10878_0 | v_10879_0;
  assign v_10878_0 = v_607_0 ? v_2566_0 : 3'h0;
  assign v_10879_0 = v_26_0 ? v_2552_0 : 3'h0;
  assign v_10880_0 = v_601_0 ? v_2545_0 : 3'h0;
  assign v_10881_0 = v_10882_0 | v_10883_0;
  assign v_10882_0 = v_607_0 ? v_2559_0 : 3'h0;
  assign v_10883_0 = v_26_0 ? v_2545_0 : 3'h0;
  assign v_10884_0 = v_601_0 ? v_2538_0 : 3'h0;
  assign v_10885_0 = v_10886_0 | v_10887_0;
  assign v_10886_0 = v_607_0 ? v_2552_0 : 3'h0;
  assign v_10887_0 = v_26_0 ? v_2538_0 : 3'h0;
  assign v_10888_0 = v_601_0 ? v_2531_0 : 3'h0;
  assign v_10889_0 = v_10890_0 | v_10891_0;
  assign v_10890_0 = v_607_0 ? v_2545_0 : 3'h0;
  assign v_10891_0 = v_26_0 ? v_2531_0 : 3'h0;
  assign v_10892_0 = v_601_0 ? v_2524_0 : 3'h0;
  assign v_10893_0 = v_10894_0 | v_10895_0;
  assign v_10894_0 = v_607_0 ? v_2538_0 : 3'h0;
  assign v_10895_0 = v_26_0 ? v_2524_0 : 3'h0;
  assign v_10896_0 = v_601_0 ? v_2517_0 : 3'h0;
  assign v_10897_0 = v_10898_0 | v_10899_0;
  assign v_10898_0 = v_607_0 ? v_2531_0 : 3'h0;
  assign v_10899_0 = v_26_0 ? v_2517_0 : 3'h0;
  assign v_10900_0 = v_601_0 ? v_2510_0 : 3'h0;
  assign v_10901_0 = v_10902_0 | v_10903_0;
  assign v_10902_0 = v_607_0 ? v_2524_0 : 3'h0;
  assign v_10903_0 = v_26_0 ? v_2510_0 : 3'h0;
  assign v_10904_0 = v_601_0 ? v_2503_0 : 3'h0;
  assign v_10905_0 = v_10906_0 | v_10907_0;
  assign v_10906_0 = v_607_0 ? v_2517_0 : 3'h0;
  assign v_10907_0 = v_26_0 ? v_2503_0 : 3'h0;
  assign v_10908_0 = v_601_0 ? v_2496_0 : 3'h0;
  assign v_10909_0 = v_10910_0 | v_10911_0;
  assign v_10910_0 = v_607_0 ? v_2510_0 : 3'h0;
  assign v_10911_0 = v_26_0 ? v_2496_0 : 3'h0;
  assign v_10912_0 = v_601_0 ? v_2489_0 : 3'h0;
  assign v_10913_0 = v_10914_0 | v_10915_0;
  assign v_10914_0 = v_607_0 ? v_2503_0 : 3'h0;
  assign v_10915_0 = v_26_0 ? v_2489_0 : 3'h0;
  assign v_10916_0 = v_601_0 ? v_2482_0 : 3'h0;
  assign v_10917_0 = v_10918_0 | v_10919_0;
  assign v_10918_0 = v_607_0 ? v_2496_0 : 3'h0;
  assign v_10919_0 = v_26_0 ? v_2482_0 : 3'h0;
  assign v_10920_0 = v_601_0 ? v_2475_0 : 3'h0;
  assign v_10921_0 = v_10922_0 | v_10923_0;
  assign v_10922_0 = v_607_0 ? v_2489_0 : 3'h0;
  assign v_10923_0 = v_26_0 ? v_2475_0 : 3'h0;
  assign v_10924_0 = v_601_0 ? v_2468_0 : 3'h0;
  assign v_10925_0 = v_10926_0 | v_10927_0;
  assign v_10926_0 = v_607_0 ? v_2482_0 : 3'h0;
  assign v_10927_0 = v_26_0 ? v_2468_0 : 3'h0;
  assign v_10928_0 = v_601_0 ? v_2461_0 : 3'h0;
  assign v_10929_0 = v_10930_0 | v_10931_0;
  assign v_10930_0 = v_607_0 ? v_2475_0 : 3'h0;
  assign v_10931_0 = v_26_0 ? v_2461_0 : 3'h0;
  assign v_10932_0 = v_601_0 ? v_2454_0 : 3'h0;
  assign v_10933_0 = v_10934_0 | v_10935_0;
  assign v_10934_0 = v_607_0 ? v_2468_0 : 3'h0;
  assign v_10935_0 = v_26_0 ? v_2454_0 : 3'h0;
  assign v_10936_0 = v_601_0 ? v_2447_0 : 3'h0;
  assign v_10937_0 = v_10938_0 | v_10939_0;
  assign v_10938_0 = v_607_0 ? v_2461_0 : 3'h0;
  assign v_10939_0 = v_26_0 ? v_2447_0 : 3'h0;
  assign v_10940_0 = v_601_0 ? v_2440_0 : 3'h0;
  assign v_10941_0 = v_10942_0 | v_10943_0;
  assign v_10942_0 = v_607_0 ? v_2454_0 : 3'h0;
  assign v_10943_0 = v_26_0 ? v_2440_0 : 3'h0;
  assign v_10944_0 = v_601_0 ? v_2433_0 : 3'h0;
  assign v_10945_0 = v_10946_0 | v_10947_0;
  assign v_10946_0 = v_607_0 ? v_2447_0 : 3'h0;
  assign v_10947_0 = v_26_0 ? v_2433_0 : 3'h0;
  assign v_10948_0 = v_601_0 ? v_2426_0 : 3'h0;
  assign v_10949_0 = v_10950_0 | v_10951_0;
  assign v_10950_0 = v_607_0 ? v_2440_0 : 3'h0;
  assign v_10951_0 = v_26_0 ? v_2426_0 : 3'h0;
  assign v_10952_0 = v_601_0 ? v_2419_0 : 3'h0;
  assign v_10953_0 = v_10954_0 | v_10955_0;
  assign v_10954_0 = v_607_0 ? v_2433_0 : 3'h0;
  assign v_10955_0 = v_26_0 ? v_2419_0 : 3'h0;
  assign v_10956_0 = v_601_0 ? v_2412_0 : 3'h0;
  assign v_10957_0 = v_10958_0 | v_10959_0;
  assign v_10958_0 = v_607_0 ? v_2426_0 : 3'h0;
  assign v_10959_0 = v_26_0 ? v_2412_0 : 3'h0;
  assign v_10960_0 = v_601_0 ? v_2405_0 : 3'h0;
  assign v_10961_0 = v_10962_0 | v_10963_0;
  assign v_10962_0 = v_607_0 ? v_2419_0 : 3'h0;
  assign v_10963_0 = v_26_0 ? v_2405_0 : 3'h0;
  assign v_10964_0 = v_601_0 ? v_2398_0 : 3'h0;
  assign v_10965_0 = v_10966_0 | v_10967_0;
  assign v_10966_0 = v_607_0 ? v_2412_0 : 3'h0;
  assign v_10967_0 = v_26_0 ? v_2398_0 : 3'h0;
  assign v_10968_0 = v_601_0 ? v_2391_0 : 3'h0;
  assign v_10969_0 = v_10970_0 | v_10971_0;
  assign v_10970_0 = v_607_0 ? v_2405_0 : 3'h0;
  assign v_10971_0 = v_26_0 ? v_2391_0 : 3'h0;
  assign v_10972_0 = v_601_0 ? v_2384_0 : 3'h0;
  assign v_10973_0 = v_10974_0 | v_10975_0;
  assign v_10974_0 = v_607_0 ? v_2398_0 : 3'h0;
  assign v_10975_0 = v_26_0 ? v_2384_0 : 3'h0;
  assign v_10976_0 = v_601_0 ? v_2377_0 : 3'h0;
  assign v_10977_0 = v_10978_0 | v_10979_0;
  assign v_10978_0 = v_607_0 ? v_2391_0 : 3'h0;
  assign v_10979_0 = v_26_0 ? v_2377_0 : 3'h0;
  assign v_10980_0 = v_601_0 ? v_2370_0 : 3'h0;
  assign v_10981_0 = v_10982_0 | v_10983_0;
  assign v_10982_0 = v_607_0 ? v_2384_0 : 3'h0;
  assign v_10983_0 = v_26_0 ? v_2370_0 : 3'h0;
  assign v_10984_0 = v_601_0 ? v_2363_0 : 3'h0;
  assign v_10985_0 = v_10986_0 | v_10987_0;
  assign v_10986_0 = v_607_0 ? v_2377_0 : 3'h0;
  assign v_10987_0 = v_26_0 ? v_2363_0 : 3'h0;
  assign v_10988_0 = v_601_0 ? v_2356_0 : 3'h0;
  assign v_10989_0 = v_10990_0 | v_10991_0;
  assign v_10990_0 = v_607_0 ? v_2370_0 : 3'h0;
  assign v_10991_0 = v_26_0 ? v_2356_0 : 3'h0;
  assign v_10992_0 = v_601_0 ? v_2349_0 : 3'h0;
  assign v_10993_0 = v_10994_0 | v_10995_0;
  assign v_10994_0 = v_607_0 ? v_2363_0 : 3'h0;
  assign v_10995_0 = v_26_0 ? v_2349_0 : 3'h0;
  assign v_10996_0 = v_601_0 ? v_2342_0 : 3'h0;
  assign v_10997_0 = v_10998_0 | v_10999_0;
  assign v_10998_0 = v_607_0 ? v_2356_0 : 3'h0;
  assign v_10999_0 = v_26_0 ? v_2342_0 : 3'h0;
  assign v_11000_0 = v_601_0 ? v_2335_0 : 3'h0;
  assign v_11001_0 = v_11002_0 | v_11003_0;
  assign v_11002_0 = v_607_0 ? v_2349_0 : 3'h0;
  assign v_11003_0 = v_26_0 ? v_2335_0 : 3'h0;
  assign v_11004_0 = v_601_0 ? v_2328_0 : 3'h0;
  assign v_11005_0 = v_11006_0 | v_11007_0;
  assign v_11006_0 = v_607_0 ? v_2342_0 : 3'h0;
  assign v_11007_0 = v_26_0 ? v_2328_0 : 3'h0;
  assign v_11008_0 = v_601_0 ? v_2321_0 : 3'h0;
  assign v_11009_0 = v_11010_0 | v_11011_0;
  assign v_11010_0 = v_607_0 ? v_2335_0 : 3'h0;
  assign v_11011_0 = v_26_0 ? v_2321_0 : 3'h0;
  assign v_11012_0 = v_601_0 ? v_2314_0 : 3'h0;
  assign v_11013_0 = v_11014_0 | v_11015_0;
  assign v_11014_0 = v_607_0 ? v_2328_0 : 3'h0;
  assign v_11015_0 = v_26_0 ? v_2314_0 : 3'h0;
  assign v_11016_0 = v_601_0 ? v_2307_0 : 3'h0;
  assign v_11017_0 = v_11018_0 | v_11019_0;
  assign v_11018_0 = v_607_0 ? v_2321_0 : 3'h0;
  assign v_11019_0 = v_26_0 ? v_2307_0 : 3'h0;
  assign v_11020_0 = v_601_0 ? v_2300_0 : 3'h0;
  assign v_11021_0 = v_11022_0 | v_11023_0;
  assign v_11022_0 = v_607_0 ? v_2314_0 : 3'h0;
  assign v_11023_0 = v_26_0 ? v_2300_0 : 3'h0;
  assign v_11024_0 = v_601_0 ? v_2293_0 : 3'h0;
  assign v_11025_0 = v_11026_0 | v_11027_0;
  assign v_11026_0 = v_607_0 ? v_2307_0 : 3'h0;
  assign v_11027_0 = v_26_0 ? v_2293_0 : 3'h0;
  assign v_11028_0 = v_601_0 ? v_2286_0 : 3'h0;
  assign v_11029_0 = v_11030_0 | v_11031_0;
  assign v_11030_0 = v_607_0 ? v_2300_0 : 3'h0;
  assign v_11031_0 = v_26_0 ? v_2286_0 : 3'h0;
  assign v_11032_0 = v_601_0 ? v_2279_0 : 3'h0;
  assign v_11033_0 = v_11034_0 | v_11035_0;
  assign v_11034_0 = v_607_0 ? v_2293_0 : 3'h0;
  assign v_11035_0 = v_26_0 ? v_2279_0 : 3'h0;
  assign v_11036_0 = v_601_0 ? v_2272_0 : 3'h0;
  assign v_11037_0 = v_11038_0 | v_11039_0;
  assign v_11038_0 = v_607_0 ? v_2286_0 : 3'h0;
  assign v_11039_0 = v_26_0 ? v_2272_0 : 3'h0;
  assign v_11040_0 = v_601_0 ? v_2265_0 : 3'h0;
  assign v_11041_0 = v_11042_0 | v_11043_0;
  assign v_11042_0 = v_607_0 ? v_2279_0 : 3'h0;
  assign v_11043_0 = v_26_0 ? v_2265_0 : 3'h0;
  assign v_11044_0 = v_601_0 ? v_2258_0 : 3'h0;
  assign v_11045_0 = v_11046_0 | v_11047_0;
  assign v_11046_0 = v_607_0 ? v_2272_0 : 3'h0;
  assign v_11047_0 = v_26_0 ? v_2258_0 : 3'h0;
  assign v_11048_0 = v_601_0 ? v_2251_0 : 3'h0;
  assign v_11049_0 = v_11050_0 | v_11051_0;
  assign v_11050_0 = v_607_0 ? v_2265_0 : 3'h0;
  assign v_11051_0 = v_26_0 ? v_2251_0 : 3'h0;
  assign v_11052_0 = v_601_0 ? v_2244_0 : 3'h0;
  assign v_11053_0 = v_11054_0 | v_11055_0;
  assign v_11054_0 = v_607_0 ? v_2258_0 : 3'h0;
  assign v_11055_0 = v_26_0 ? v_2244_0 : 3'h0;
  assign v_11056_0 = v_601_0 ? v_2237_0 : 3'h0;
  assign v_11057_0 = v_11058_0 | v_11059_0;
  assign v_11058_0 = v_607_0 ? v_2251_0 : 3'h0;
  assign v_11059_0 = v_26_0 ? v_2237_0 : 3'h0;
  assign v_11060_0 = v_601_0 ? v_2230_0 : 3'h0;
  assign v_11061_0 = v_11062_0 | v_11063_0;
  assign v_11062_0 = v_607_0 ? v_2244_0 : 3'h0;
  assign v_11063_0 = v_26_0 ? v_2230_0 : 3'h0;
  assign v_11064_0 = v_601_0 ? v_2223_0 : 3'h0;
  assign v_11065_0 = v_11066_0 | v_11067_0;
  assign v_11066_0 = v_607_0 ? v_2237_0 : 3'h0;
  assign v_11067_0 = v_26_0 ? v_2223_0 : 3'h0;
  assign v_11068_0 = v_601_0 ? v_2216_0 : 3'h0;
  assign v_11069_0 = v_11070_0 | v_11071_0;
  assign v_11070_0 = v_607_0 ? v_2230_0 : 3'h0;
  assign v_11071_0 = v_26_0 ? v_2216_0 : 3'h0;
  assign v_11072_0 = v_601_0 ? v_2209_0 : 3'h0;
  assign v_11073_0 = v_11074_0 | v_11075_0;
  assign v_11074_0 = v_607_0 ? v_2223_0 : 3'h0;
  assign v_11075_0 = v_26_0 ? v_2209_0 : 3'h0;
  assign v_11076_0 = v_601_0 ? v_2202_0 : 3'h0;
  assign v_11077_0 = v_11078_0 | v_11079_0;
  assign v_11078_0 = v_607_0 ? v_2216_0 : 3'h0;
  assign v_11079_0 = v_26_0 ? v_2202_0 : 3'h0;
  assign v_11080_0 = v_601_0 ? v_2195_0 : 3'h0;
  assign v_11081_0 = v_11082_0 | v_11083_0;
  assign v_11082_0 = v_607_0 ? v_2209_0 : 3'h0;
  assign v_11083_0 = v_26_0 ? v_2195_0 : 3'h0;
  assign v_11084_0 = v_601_0 ? v_2188_0 : 3'h0;
  assign v_11085_0 = v_11086_0 | v_11087_0;
  assign v_11086_0 = v_607_0 ? v_2202_0 : 3'h0;
  assign v_11087_0 = v_26_0 ? v_2188_0 : 3'h0;
  assign v_11088_0 = v_601_0 ? v_2181_0 : 3'h0;
  assign v_11089_0 = v_11090_0 | v_11091_0;
  assign v_11090_0 = v_607_0 ? v_2195_0 : 3'h0;
  assign v_11091_0 = v_26_0 ? v_2181_0 : 3'h0;
  assign v_11092_0 = v_601_0 ? v_2174_0 : 3'h0;
  assign v_11093_0 = v_11094_0 | v_11095_0;
  assign v_11094_0 = v_607_0 ? v_2188_0 : 3'h0;
  assign v_11095_0 = v_26_0 ? v_2174_0 : 3'h0;
  assign v_11096_0 = v_601_0 ? v_2167_0 : 3'h0;
  assign v_11097_0 = v_11098_0 | v_11099_0;
  assign v_11098_0 = v_607_0 ? v_2181_0 : 3'h0;
  assign v_11099_0 = v_26_0 ? v_2167_0 : 3'h0;
  assign v_11100_0 = v_601_0 ? v_2160_0 : 3'h0;
  assign v_11101_0 = v_11102_0 | v_11103_0;
  assign v_11102_0 = v_607_0 ? v_2174_0 : 3'h0;
  assign v_11103_0 = v_26_0 ? v_2160_0 : 3'h0;
  assign v_11104_0 = v_601_0 ? v_2153_0 : 3'h0;
  assign v_11105_0 = v_11106_0 | v_11107_0;
  assign v_11106_0 = v_607_0 ? v_2167_0 : 3'h0;
  assign v_11107_0 = v_26_0 ? v_2153_0 : 3'h0;
  assign v_11108_0 = v_601_0 ? v_2146_0 : 3'h0;
  assign v_11109_0 = v_11110_0 | v_11111_0;
  assign v_11110_0 = v_607_0 ? v_2160_0 : 3'h0;
  assign v_11111_0 = v_26_0 ? v_2146_0 : 3'h0;
  assign v_11112_0 = v_601_0 ? v_2139_0 : 3'h0;
  assign v_11113_0 = v_11114_0 | v_11115_0;
  assign v_11114_0 = v_607_0 ? v_2153_0 : 3'h0;
  assign v_11115_0 = v_26_0 ? v_2139_0 : 3'h0;
  assign v_11116_0 = v_601_0 ? v_2132_0 : 3'h0;
  assign v_11117_0 = v_11118_0 | v_11119_0;
  assign v_11118_0 = v_607_0 ? v_2146_0 : 3'h0;
  assign v_11119_0 = v_26_0 ? v_2132_0 : 3'h0;
  assign v_11120_0 = v_601_0 ? v_2125_0 : 3'h0;
  assign v_11121_0 = v_11122_0 | v_11123_0;
  assign v_11122_0 = v_607_0 ? v_2139_0 : 3'h0;
  assign v_11123_0 = v_26_0 ? v_2125_0 : 3'h0;
  assign v_11124_0 = v_601_0 ? v_2118_0 : 3'h0;
  assign v_11125_0 = v_11126_0 | v_11127_0;
  assign v_11126_0 = v_607_0 ? v_2132_0 : 3'h0;
  assign v_11127_0 = v_26_0 ? v_2118_0 : 3'h0;
  assign v_11128_0 = v_601_0 ? v_2111_0 : 3'h0;
  assign v_11129_0 = v_11130_0 | v_11131_0;
  assign v_11130_0 = v_607_0 ? v_2125_0 : 3'h0;
  assign v_11131_0 = v_26_0 ? v_2111_0 : 3'h0;
  assign v_11132_0 = v_601_0 ? v_2104_0 : 3'h0;
  assign v_11133_0 = v_11134_0 | v_11135_0;
  assign v_11134_0 = v_607_0 ? v_2118_0 : 3'h0;
  assign v_11135_0 = v_26_0 ? v_2104_0 : 3'h0;
  assign v_11136_0 = v_601_0 ? v_2097_0 : 3'h0;
  assign v_11137_0 = v_11138_0 | v_11139_0;
  assign v_11138_0 = v_607_0 ? v_2111_0 : 3'h0;
  assign v_11139_0 = v_26_0 ? v_2097_0 : 3'h0;
  assign v_11140_0 = v_601_0 ? v_2090_0 : 3'h0;
  assign v_11141_0 = v_11142_0 | v_11143_0;
  assign v_11142_0 = v_607_0 ? v_2104_0 : 3'h0;
  assign v_11143_0 = v_26_0 ? v_2090_0 : 3'h0;
  assign v_11144_0 = v_601_0 ? v_2083_0 : 3'h0;
  assign v_11145_0 = v_11146_0 | v_11147_0;
  assign v_11146_0 = v_607_0 ? v_2097_0 : 3'h0;
  assign v_11147_0 = v_26_0 ? v_2083_0 : 3'h0;
  assign v_11148_0 = v_601_0 ? v_2076_0 : 3'h0;
  assign v_11149_0 = v_11150_0 | v_11151_0;
  assign v_11150_0 = v_607_0 ? v_2090_0 : 3'h0;
  assign v_11151_0 = v_26_0 ? v_2076_0 : 3'h0;
  assign v_11152_0 = v_601_0 ? v_2069_0 : 3'h0;
  assign v_11153_0 = v_11154_0 | v_11155_0;
  assign v_11154_0 = v_607_0 ? v_2083_0 : 3'h0;
  assign v_11155_0 = v_26_0 ? v_2069_0 : 3'h0;
  assign v_11156_0 = v_601_0 ? v_2062_0 : 3'h0;
  assign v_11157_0 = v_11158_0 | v_11159_0;
  assign v_11158_0 = v_607_0 ? v_2076_0 : 3'h0;
  assign v_11159_0 = v_26_0 ? v_2062_0 : 3'h0;
  assign v_11160_0 = v_601_0 ? v_2055_0 : 3'h0;
  assign v_11161_0 = v_11162_0 | v_11163_0;
  assign v_11162_0 = v_607_0 ? v_2069_0 : 3'h0;
  assign v_11163_0 = v_26_0 ? v_2055_0 : 3'h0;
  assign v_11164_0 = v_601_0 ? v_2048_0 : 3'h0;
  assign v_11165_0 = v_11166_0 | v_11167_0;
  assign v_11166_0 = v_607_0 ? v_2062_0 : 3'h0;
  assign v_11167_0 = v_26_0 ? v_2048_0 : 3'h0;
  assign v_11168_0 = v_601_0 ? v_2041_0 : 3'h0;
  assign v_11169_0 = v_11170_0 | v_11171_0;
  assign v_11170_0 = v_607_0 ? v_2055_0 : 3'h0;
  assign v_11171_0 = v_26_0 ? v_2041_0 : 3'h0;
  assign v_11172_0 = v_601_0 ? v_2034_0 : 3'h0;
  assign v_11173_0 = v_11174_0 | v_11175_0;
  assign v_11174_0 = v_607_0 ? v_2048_0 : 3'h0;
  assign v_11175_0 = v_26_0 ? v_2034_0 : 3'h0;
  assign v_11176_0 = v_601_0 ? v_2027_0 : 3'h0;
  assign v_11177_0 = v_11178_0 | v_11179_0;
  assign v_11178_0 = v_607_0 ? v_2041_0 : 3'h0;
  assign v_11179_0 = v_26_0 ? v_2027_0 : 3'h0;
  assign v_11180_0 = v_601_0 ? v_2020_0 : 3'h0;
  assign v_11181_0 = v_11182_0 | v_11183_0;
  assign v_11182_0 = v_607_0 ? v_2034_0 : 3'h0;
  assign v_11183_0 = v_26_0 ? v_2020_0 : 3'h0;
  assign v_11184_0 = v_601_0 ? v_2013_0 : 3'h0;
  assign v_11185_0 = v_11186_0 | v_11187_0;
  assign v_11186_0 = v_607_0 ? v_2027_0 : 3'h0;
  assign v_11187_0 = v_26_0 ? v_2013_0 : 3'h0;
  assign v_11188_0 = v_601_0 ? v_2006_0 : 3'h0;
  assign v_11189_0 = v_11190_0 | v_11191_0;
  assign v_11190_0 = v_607_0 ? v_2020_0 : 3'h0;
  assign v_11191_0 = v_26_0 ? v_2006_0 : 3'h0;
  assign v_11192_0 = v_601_0 ? v_1999_0 : 3'h0;
  assign v_11193_0 = v_11194_0 | v_11195_0;
  assign v_11194_0 = v_607_0 ? v_2013_0 : 3'h0;
  assign v_11195_0 = v_26_0 ? v_1999_0 : 3'h0;
  assign v_11196_0 = v_601_0 ? v_1992_0 : 3'h0;
  assign v_11197_0 = v_11198_0 | v_11199_0;
  assign v_11198_0 = v_607_0 ? v_2006_0 : 3'h0;
  assign v_11199_0 = v_26_0 ? v_1992_0 : 3'h0;
  assign v_11200_0 = v_601_0 ? v_1985_0 : 3'h0;
  assign v_11201_0 = v_11202_0 | v_11203_0;
  assign v_11202_0 = v_607_0 ? v_1999_0 : 3'h0;
  assign v_11203_0 = v_26_0 ? v_1985_0 : 3'h0;
  assign v_11204_0 = v_601_0 ? v_1978_0 : 3'h0;
  assign v_11205_0 = v_11206_0 | v_11207_0;
  assign v_11206_0 = v_607_0 ? v_1992_0 : 3'h0;
  assign v_11207_0 = v_26_0 ? v_1978_0 : 3'h0;
  assign v_11208_0 = v_601_0 ? v_1971_0 : 3'h0;
  assign v_11209_0 = v_11210_0 | v_11211_0;
  assign v_11210_0 = v_607_0 ? v_1985_0 : 3'h0;
  assign v_11211_0 = v_26_0 ? v_1971_0 : 3'h0;
  assign v_11212_0 = v_601_0 ? v_1964_0 : 3'h0;
  assign v_11213_0 = v_11214_0 | v_11215_0;
  assign v_11214_0 = v_607_0 ? v_1978_0 : 3'h0;
  assign v_11215_0 = v_26_0 ? v_1964_0 : 3'h0;
  assign v_11216_0 = v_601_0 ? v_1957_0 : 3'h0;
  assign v_11217_0 = v_11218_0 | v_11219_0;
  assign v_11218_0 = v_607_0 ? v_1971_0 : 3'h0;
  assign v_11219_0 = v_26_0 ? v_1957_0 : 3'h0;
  assign v_11220_0 = v_601_0 ? v_1950_0 : 3'h0;
  assign v_11221_0 = v_11222_0 | v_11223_0;
  assign v_11222_0 = v_607_0 ? v_1964_0 : 3'h0;
  assign v_11223_0 = v_26_0 ? v_1950_0 : 3'h0;
  assign v_11224_0 = v_601_0 ? v_1943_0 : 3'h0;
  assign v_11225_0 = v_11226_0 | v_11227_0;
  assign v_11226_0 = v_607_0 ? v_1957_0 : 3'h0;
  assign v_11227_0 = v_26_0 ? v_1943_0 : 3'h0;
  assign v_11228_0 = v_601_0 ? v_1936_0 : 3'h0;
  assign v_11229_0 = v_11230_0 | v_11231_0;
  assign v_11230_0 = v_607_0 ? v_1950_0 : 3'h0;
  assign v_11231_0 = v_26_0 ? v_1936_0 : 3'h0;
  assign v_11232_0 = v_601_0 ? v_1929_0 : 3'h0;
  assign v_11233_0 = v_11234_0 | v_11235_0;
  assign v_11234_0 = v_607_0 ? v_1943_0 : 3'h0;
  assign v_11235_0 = v_26_0 ? v_1929_0 : 3'h0;
  assign v_11236_0 = v_601_0 ? v_1922_0 : 3'h0;
  assign v_11237_0 = v_11238_0 | v_11239_0;
  assign v_11238_0 = v_607_0 ? v_1936_0 : 3'h0;
  assign v_11239_0 = v_26_0 ? v_1922_0 : 3'h0;
  assign v_11240_0 = v_601_0 ? v_1915_0 : 3'h0;
  assign v_11241_0 = v_11242_0 | v_11243_0;
  assign v_11242_0 = v_607_0 ? v_1929_0 : 3'h0;
  assign v_11243_0 = v_26_0 ? v_1915_0 : 3'h0;
  assign v_11244_0 = v_601_0 ? v_1908_0 : 3'h0;
  assign v_11245_0 = v_11246_0 | v_11247_0;
  assign v_11246_0 = v_607_0 ? v_1922_0 : 3'h0;
  assign v_11247_0 = v_26_0 ? v_1908_0 : 3'h0;
  assign v_11248_0 = v_601_0 ? v_1901_0 : 3'h0;
  assign v_11249_0 = v_11250_0 | v_11251_0;
  assign v_11250_0 = v_607_0 ? v_1915_0 : 3'h0;
  assign v_11251_0 = v_26_0 ? v_1901_0 : 3'h0;
  assign v_11252_0 = v_601_0 ? v_1894_0 : 3'h0;
  assign v_11253_0 = v_11254_0 | v_11255_0;
  assign v_11254_0 = v_607_0 ? v_1908_0 : 3'h0;
  assign v_11255_0 = v_26_0 ? v_1894_0 : 3'h0;
  assign v_11256_0 = v_601_0 ? v_1887_0 : 3'h0;
  assign v_11257_0 = v_11258_0 | v_11259_0;
  assign v_11258_0 = v_607_0 ? v_1901_0 : 3'h0;
  assign v_11259_0 = v_26_0 ? v_1887_0 : 3'h0;
  assign v_11260_0 = v_601_0 ? v_1880_0 : 3'h0;
  assign v_11261_0 = v_11262_0 | v_11263_0;
  assign v_11262_0 = v_607_0 ? v_1894_0 : 3'h0;
  assign v_11263_0 = v_26_0 ? v_1880_0 : 3'h0;
  assign v_11264_0 = v_601_0 ? v_1873_0 : 3'h0;
  assign v_11265_0 = v_11266_0 | v_11267_0;
  assign v_11266_0 = v_607_0 ? v_1887_0 : 3'h0;
  assign v_11267_0 = v_26_0 ? v_1873_0 : 3'h0;
  assign v_11268_0 = v_601_0 ? v_1866_0 : 3'h0;
  assign v_11269_0 = v_11270_0 | v_11271_0;
  assign v_11270_0 = v_607_0 ? v_1880_0 : 3'h0;
  assign v_11271_0 = v_26_0 ? v_1866_0 : 3'h0;
  assign v_11272_0 = v_601_0 ? v_1859_0 : 3'h0;
  assign v_11273_0 = v_11274_0 | v_11275_0;
  assign v_11274_0 = v_607_0 ? v_1873_0 : 3'h0;
  assign v_11275_0 = v_26_0 ? v_1859_0 : 3'h0;
  assign v_11276_0 = v_601_0 ? v_1852_0 : 3'h0;
  assign v_11277_0 = v_11278_0 | v_11279_0;
  assign v_11278_0 = v_607_0 ? v_1866_0 : 3'h0;
  assign v_11279_0 = v_26_0 ? v_1852_0 : 3'h0;
  assign v_11280_0 = v_601_0 ? v_1845_0 : 3'h0;
  assign v_11281_0 = v_11282_0 | v_11283_0;
  assign v_11282_0 = v_607_0 ? v_1859_0 : 3'h0;
  assign v_11283_0 = v_26_0 ? v_1845_0 : 3'h0;
  assign v_11284_0 = v_601_0 ? v_1838_0 : 3'h0;
  assign v_11285_0 = v_11286_0 | v_11287_0;
  assign v_11286_0 = v_607_0 ? v_1852_0 : 3'h0;
  assign v_11287_0 = v_26_0 ? v_1838_0 : 3'h0;
  assign v_11288_0 = v_601_0 ? v_1831_0 : 3'h0;
  assign v_11289_0 = v_11290_0 | v_11291_0;
  assign v_11290_0 = v_607_0 ? v_1845_0 : 3'h0;
  assign v_11291_0 = v_26_0 ? v_1831_0 : 3'h0;
  assign v_11292_0 = v_601_0 ? v_1824_0 : 3'h0;
  assign v_11293_0 = v_11294_0 | v_11295_0;
  assign v_11294_0 = v_607_0 ? v_1838_0 : 3'h0;
  assign v_11295_0 = v_26_0 ? v_1824_0 : 3'h0;
  assign v_11296_0 = v_601_0 ? v_1817_0 : 3'h0;
  assign v_11297_0 = v_11298_0 | v_11299_0;
  assign v_11298_0 = v_607_0 ? v_1831_0 : 3'h0;
  assign v_11299_0 = v_26_0 ? v_1817_0 : 3'h0;
  assign v_11300_0 = v_601_0 ? v_1810_0 : 3'h0;
  assign v_11301_0 = v_11302_0 | v_11303_0;
  assign v_11302_0 = v_607_0 ? v_1824_0 : 3'h0;
  assign v_11303_0 = v_26_0 ? v_1810_0 : 3'h0;
  assign v_11304_0 = v_601_0 ? v_1803_0 : 3'h0;
  assign v_11305_0 = v_11306_0 | v_11307_0;
  assign v_11306_0 = v_607_0 ? v_1817_0 : 3'h0;
  assign v_11307_0 = v_26_0 ? v_1803_0 : 3'h0;
  assign v_11308_0 = v_601_0 ? v_1796_0 : 3'h0;
  assign v_11309_0 = v_11310_0 | v_11311_0;
  assign v_11310_0 = v_607_0 ? v_1810_0 : 3'h0;
  assign v_11311_0 = v_26_0 ? v_1796_0 : 3'h0;
  assign v_11312_0 = v_601_0 ? v_1789_0 : 3'h0;
  assign v_11313_0 = v_11314_0 | v_11315_0;
  assign v_11314_0 = v_607_0 ? v_1803_0 : 3'h0;
  assign v_11315_0 = v_26_0 ? v_1789_0 : 3'h0;
  assign v_11316_0 = v_601_0 ? v_1782_0 : 3'h0;
  assign v_11317_0 = v_11318_0 | v_11319_0;
  assign v_11318_0 = v_607_0 ? v_1796_0 : 3'h0;
  assign v_11319_0 = v_26_0 ? v_1782_0 : 3'h0;
  assign v_11320_0 = v_601_0 ? v_1775_0 : 3'h0;
  assign v_11321_0 = v_11322_0 | v_11323_0;
  assign v_11322_0 = v_607_0 ? v_1789_0 : 3'h0;
  assign v_11323_0 = v_26_0 ? v_1775_0 : 3'h0;
  assign v_11324_0 = v_601_0 ? v_1768_0 : 3'h0;
  assign v_11325_0 = v_11326_0 | v_11327_0;
  assign v_11326_0 = v_607_0 ? v_1782_0 : 3'h0;
  assign v_11327_0 = v_26_0 ? v_1768_0 : 3'h0;
  assign v_11328_0 = v_601_0 ? v_1761_0 : 3'h0;
  assign v_11329_0 = v_11330_0 | v_11331_0;
  assign v_11330_0 = v_607_0 ? v_1775_0 : 3'h0;
  assign v_11331_0 = v_26_0 ? v_1761_0 : 3'h0;
  assign v_11332_0 = v_601_0 ? v_1754_0 : 3'h0;
  assign v_11333_0 = v_11334_0 | v_11335_0;
  assign v_11334_0 = v_607_0 ? v_1768_0 : 3'h0;
  assign v_11335_0 = v_26_0 ? v_1754_0 : 3'h0;
  assign v_11336_0 = v_601_0 ? v_1747_0 : 3'h0;
  assign v_11337_0 = v_11338_0 | v_11339_0;
  assign v_11338_0 = v_607_0 ? v_1761_0 : 3'h0;
  assign v_11339_0 = v_26_0 ? v_1747_0 : 3'h0;
  assign v_11340_0 = v_601_0 ? v_1740_0 : 3'h0;
  assign v_11341_0 = v_11342_0 | v_11343_0;
  assign v_11342_0 = v_607_0 ? v_1754_0 : 3'h0;
  assign v_11343_0 = v_26_0 ? v_1740_0 : 3'h0;
  assign v_11344_0 = v_601_0 ? v_1733_0 : 3'h0;
  assign v_11345_0 = v_11346_0 | v_11347_0;
  assign v_11346_0 = v_607_0 ? v_1747_0 : 3'h0;
  assign v_11347_0 = v_26_0 ? v_1733_0 : 3'h0;
  assign v_11348_0 = v_601_0 ? v_1726_0 : 3'h0;
  assign v_11349_0 = v_11350_0 | v_11351_0;
  assign v_11350_0 = v_607_0 ? v_1740_0 : 3'h0;
  assign v_11351_0 = v_26_0 ? v_1726_0 : 3'h0;
  assign v_11352_0 = v_601_0 ? v_1719_0 : 3'h0;
  assign v_11353_0 = v_11354_0 | v_11355_0;
  assign v_11354_0 = v_607_0 ? v_1733_0 : 3'h0;
  assign v_11355_0 = v_26_0 ? v_1719_0 : 3'h0;
  assign v_11356_0 = v_601_0 ? v_1712_0 : 3'h0;
  assign v_11357_0 = v_11358_0 | v_11359_0;
  assign v_11358_0 = v_607_0 ? v_1726_0 : 3'h0;
  assign v_11359_0 = v_26_0 ? v_1712_0 : 3'h0;
  assign v_11360_0 = v_601_0 ? v_1705_0 : 3'h0;
  assign v_11361_0 = v_11362_0 | v_11363_0;
  assign v_11362_0 = v_607_0 ? v_1719_0 : 3'h0;
  assign v_11363_0 = v_26_0 ? v_1705_0 : 3'h0;
  assign v_11364_0 = v_601_0 ? v_1698_0 : 3'h0;
  assign v_11365_0 = v_11366_0 | v_11367_0;
  assign v_11366_0 = v_607_0 ? v_1712_0 : 3'h0;
  assign v_11367_0 = v_26_0 ? v_1698_0 : 3'h0;
  assign v_11368_0 = v_601_0 ? v_1691_0 : 3'h0;
  assign v_11369_0 = v_11370_0 | v_11371_0;
  assign v_11370_0 = v_607_0 ? v_1705_0 : 3'h0;
  assign v_11371_0 = v_26_0 ? v_1691_0 : 3'h0;
  assign v_11372_0 = v_601_0 ? v_1684_0 : 3'h0;
  assign v_11373_0 = v_11374_0 | v_11375_0;
  assign v_11374_0 = v_607_0 ? v_1698_0 : 3'h0;
  assign v_11375_0 = v_26_0 ? v_1684_0 : 3'h0;
  assign v_11376_0 = v_601_0 ? v_1677_0 : 3'h0;
  assign v_11377_0 = v_11378_0 | v_11379_0;
  assign v_11378_0 = v_607_0 ? v_1691_0 : 3'h0;
  assign v_11379_0 = v_26_0 ? v_1677_0 : 3'h0;
  assign v_11380_0 = v_601_0 ? v_1670_0 : 3'h0;
  assign v_11381_0 = v_11382_0 | v_11383_0;
  assign v_11382_0 = v_607_0 ? v_1684_0 : 3'h0;
  assign v_11383_0 = v_26_0 ? v_1670_0 : 3'h0;
  assign v_11384_0 = v_601_0 ? v_1663_0 : 3'h0;
  assign v_11385_0 = v_11386_0 | v_11387_0;
  assign v_11386_0 = v_607_0 ? v_1677_0 : 3'h0;
  assign v_11387_0 = v_26_0 ? v_1663_0 : 3'h0;
  assign v_11388_0 = v_601_0 ? v_1656_0 : 3'h0;
  assign v_11389_0 = v_11390_0 | v_11391_0;
  assign v_11390_0 = v_607_0 ? v_1670_0 : 3'h0;
  assign v_11391_0 = v_26_0 ? v_1656_0 : 3'h0;
  assign v_11392_0 = v_601_0 ? v_1649_0 : 3'h0;
  assign v_11393_0 = v_11394_0 | v_11395_0;
  assign v_11394_0 = v_607_0 ? v_1663_0 : 3'h0;
  assign v_11395_0 = v_26_0 ? v_1649_0 : 3'h0;
  assign v_11396_0 = v_601_0 ? v_1642_0 : 3'h0;
  assign v_11397_0 = v_11398_0 | v_11399_0;
  assign v_11398_0 = v_607_0 ? v_1656_0 : 3'h0;
  assign v_11399_0 = v_26_0 ? v_1642_0 : 3'h0;
  assign v_11400_0 = v_601_0 ? v_1635_0 : 3'h0;
  assign v_11401_0 = v_11402_0 | v_11403_0;
  assign v_11402_0 = v_607_0 ? v_1649_0 : 3'h0;
  assign v_11403_0 = v_26_0 ? v_1635_0 : 3'h0;
  assign v_11404_0 = v_601_0 ? v_1628_0 : 3'h0;
  assign v_11405_0 = v_11406_0 | v_11407_0;
  assign v_11406_0 = v_607_0 ? v_1642_0 : 3'h0;
  assign v_11407_0 = v_26_0 ? v_1628_0 : 3'h0;
  assign v_11408_0 = v_601_0 ? v_1621_0 : 3'h0;
  assign v_11409_0 = v_11410_0 | v_11411_0;
  assign v_11410_0 = v_607_0 ? v_1635_0 : 3'h0;
  assign v_11411_0 = v_26_0 ? v_1621_0 : 3'h0;
  assign v_11412_0 = v_601_0 ? v_1614_0 : 3'h0;
  assign v_11413_0 = v_11414_0 | v_11415_0;
  assign v_11414_0 = v_607_0 ? v_1628_0 : 3'h0;
  assign v_11415_0 = v_26_0 ? v_1614_0 : 3'h0;
  assign v_11416_0 = v_601_0 ? v_1607_0 : 3'h0;
  assign v_11417_0 = v_11418_0 | v_11419_0;
  assign v_11418_0 = v_607_0 ? v_1621_0 : 3'h0;
  assign v_11419_0 = v_26_0 ? v_1607_0 : 3'h0;
  assign v_11420_0 = v_601_0 ? v_1600_0 : 3'h0;
  assign v_11421_0 = v_11422_0 | v_11423_0;
  assign v_11422_0 = v_607_0 ? v_1614_0 : 3'h0;
  assign v_11423_0 = v_26_0 ? v_1600_0 : 3'h0;
  assign v_11424_0 = v_601_0 ? v_1593_0 : 3'h0;
  assign v_11425_0 = v_11426_0 | v_11427_0;
  assign v_11426_0 = v_607_0 ? v_1607_0 : 3'h0;
  assign v_11427_0 = v_26_0 ? v_1593_0 : 3'h0;
  assign v_11428_0 = v_601_0 ? v_1586_0 : 3'h0;
  assign v_11429_0 = v_11430_0 | v_11431_0;
  assign v_11430_0 = v_607_0 ? v_1600_0 : 3'h0;
  assign v_11431_0 = v_26_0 ? v_1586_0 : 3'h0;
  assign v_11432_0 = v_601_0 ? v_1579_0 : 3'h0;
  assign v_11433_0 = v_11434_0 | v_11435_0;
  assign v_11434_0 = v_607_0 ? v_1593_0 : 3'h0;
  assign v_11435_0 = v_26_0 ? v_1579_0 : 3'h0;
  assign v_11436_0 = v_601_0 ? v_1572_0 : 3'h0;
  assign v_11437_0 = v_11438_0 | v_11439_0;
  assign v_11438_0 = v_607_0 ? v_1586_0 : 3'h0;
  assign v_11439_0 = v_26_0 ? v_1572_0 : 3'h0;
  assign v_11440_0 = v_601_0 ? v_1565_0 : 3'h0;
  assign v_11441_0 = v_11442_0 | v_11443_0;
  assign v_11442_0 = v_607_0 ? v_1579_0 : 3'h0;
  assign v_11443_0 = v_26_0 ? v_1565_0 : 3'h0;
  assign v_11444_0 = v_601_0 ? v_1558_0 : 3'h0;
  assign v_11445_0 = v_11446_0 | v_11447_0;
  assign v_11446_0 = v_607_0 ? v_1572_0 : 3'h0;
  assign v_11447_0 = v_26_0 ? v_1558_0 : 3'h0;
  assign v_11448_0 = v_601_0 ? v_1551_0 : 3'h0;
  assign v_11449_0 = v_11450_0 | v_11451_0;
  assign v_11450_0 = v_607_0 ? v_1565_0 : 3'h0;
  assign v_11451_0 = v_26_0 ? v_1551_0 : 3'h0;
  assign v_11452_0 = v_601_0 ? v_1544_0 : 3'h0;
  assign v_11453_0 = v_11454_0 | v_11455_0;
  assign v_11454_0 = v_607_0 ? v_1558_0 : 3'h0;
  assign v_11455_0 = v_26_0 ? v_1544_0 : 3'h0;
  assign v_11456_0 = v_601_0 ? v_1537_0 : 3'h0;
  assign v_11457_0 = v_11458_0 | v_11459_0;
  assign v_11458_0 = v_607_0 ? v_1551_0 : 3'h0;
  assign v_11459_0 = v_26_0 ? v_1537_0 : 3'h0;
  assign v_11460_0 = v_601_0 ? v_1530_0 : 3'h0;
  assign v_11461_0 = v_11462_0 | v_11463_0;
  assign v_11462_0 = v_607_0 ? v_1544_0 : 3'h0;
  assign v_11463_0 = v_26_0 ? v_1530_0 : 3'h0;
  assign v_11464_0 = v_601_0 ? v_1523_0 : 3'h0;
  assign v_11465_0 = v_11466_0 | v_11467_0;
  assign v_11466_0 = v_607_0 ? v_1537_0 : 3'h0;
  assign v_11467_0 = v_26_0 ? v_1523_0 : 3'h0;
  assign v_11468_0 = v_601_0 ? v_1516_0 : 3'h0;
  assign v_11469_0 = v_11470_0 | v_11471_0;
  assign v_11470_0 = v_607_0 ? v_1530_0 : 3'h0;
  assign v_11471_0 = v_26_0 ? v_1516_0 : 3'h0;
  assign v_11472_0 = v_601_0 ? v_1509_0 : 3'h0;
  assign v_11473_0 = v_11474_0 | v_11475_0;
  assign v_11474_0 = v_607_0 ? v_1523_0 : 3'h0;
  assign v_11475_0 = v_26_0 ? v_1509_0 : 3'h0;
  assign v_11476_0 = v_601_0 ? v_1502_0 : 3'h0;
  assign v_11477_0 = v_11478_0 | v_11479_0;
  assign v_11478_0 = v_607_0 ? v_1516_0 : 3'h0;
  assign v_11479_0 = v_26_0 ? v_1502_0 : 3'h0;
  assign v_11480_0 = v_601_0 ? v_1495_0 : 3'h0;
  assign v_11481_0 = v_11482_0 | v_11483_0;
  assign v_11482_0 = v_607_0 ? v_1509_0 : 3'h0;
  assign v_11483_0 = v_26_0 ? v_1495_0 : 3'h0;
  assign v_11484_0 = v_601_0 ? v_1488_0 : 3'h0;
  assign v_11485_0 = v_11486_0 | v_11487_0;
  assign v_11486_0 = v_607_0 ? v_1502_0 : 3'h0;
  assign v_11487_0 = v_26_0 ? v_1488_0 : 3'h0;
  assign v_11488_0 = v_601_0 ? v_1481_0 : 3'h0;
  assign v_11489_0 = v_11490_0 | v_11491_0;
  assign v_11490_0 = v_607_0 ? v_1495_0 : 3'h0;
  assign v_11491_0 = v_26_0 ? v_1481_0 : 3'h0;
  assign v_11492_0 = v_601_0 ? v_1474_0 : 3'h0;
  assign v_11493_0 = v_11494_0 | v_11495_0;
  assign v_11494_0 = v_607_0 ? v_1488_0 : 3'h0;
  assign v_11495_0 = v_26_0 ? v_1474_0 : 3'h0;
  assign v_11496_0 = v_601_0 ? v_1467_0 : 3'h0;
  assign v_11497_0 = v_11498_0 | v_11499_0;
  assign v_11498_0 = v_607_0 ? v_1481_0 : 3'h0;
  assign v_11499_0 = v_26_0 ? v_1467_0 : 3'h0;
  assign v_11500_0 = v_601_0 ? v_1460_0 : 3'h0;
  assign v_11501_0 = v_11502_0 | v_11503_0;
  assign v_11502_0 = v_607_0 ? v_1474_0 : 3'h0;
  assign v_11503_0 = v_26_0 ? v_1460_0 : 3'h0;
  assign v_11504_0 = v_601_0 ? v_1453_0 : 3'h0;
  assign v_11505_0 = v_11506_0 | v_11507_0;
  assign v_11506_0 = v_607_0 ? v_1467_0 : 3'h0;
  assign v_11507_0 = v_26_0 ? v_1453_0 : 3'h0;
  assign v_11508_0 = v_601_0 ? v_1446_0 : 3'h0;
  assign v_11509_0 = v_11510_0 | v_11511_0;
  assign v_11510_0 = v_607_0 ? v_1460_0 : 3'h0;
  assign v_11511_0 = v_26_0 ? v_1446_0 : 3'h0;
  assign v_11512_0 = v_601_0 ? v_1439_0 : 3'h0;
  assign v_11513_0 = v_11514_0 | v_11515_0;
  assign v_11514_0 = v_607_0 ? v_1453_0 : 3'h0;
  assign v_11515_0 = v_26_0 ? v_1439_0 : 3'h0;
  assign v_11516_0 = v_601_0 ? v_1432_0 : 3'h0;
  assign v_11517_0 = v_11518_0 | v_11519_0;
  assign v_11518_0 = v_607_0 ? v_1446_0 : 3'h0;
  assign v_11519_0 = v_26_0 ? v_1432_0 : 3'h0;
  assign v_11520_0 = v_601_0 ? v_1425_0 : 3'h0;
  assign v_11521_0 = v_11522_0 | v_11523_0;
  assign v_11522_0 = v_607_0 ? v_1439_0 : 3'h0;
  assign v_11523_0 = v_26_0 ? v_1425_0 : 3'h0;
  assign v_11524_0 = v_601_0 ? v_1418_0 : 3'h0;
  assign v_11525_0 = v_11526_0 | v_11527_0;
  assign v_11526_0 = v_607_0 ? v_1432_0 : 3'h0;
  assign v_11527_0 = v_26_0 ? v_1418_0 : 3'h0;
  assign v_11528_0 = v_601_0 ? v_1411_0 : 3'h0;
  assign v_11529_0 = v_11530_0 | v_11531_0;
  assign v_11530_0 = v_607_0 ? v_1425_0 : 3'h0;
  assign v_11531_0 = v_26_0 ? v_1411_0 : 3'h0;
  assign v_11532_0 = v_601_0 ? v_1404_0 : 3'h0;
  assign v_11533_0 = v_11534_0 | v_11535_0;
  assign v_11534_0 = v_607_0 ? v_1418_0 : 3'h0;
  assign v_11535_0 = v_26_0 ? v_1404_0 : 3'h0;
  assign v_11536_0 = v_601_0 ? v_1397_0 : 3'h0;
  assign v_11537_0 = v_11538_0 | v_11539_0;
  assign v_11538_0 = v_607_0 ? v_1411_0 : 3'h0;
  assign v_11539_0 = v_26_0 ? v_1397_0 : 3'h0;
  assign v_11540_0 = v_601_0 ? v_1390_0 : 3'h0;
  assign v_11541_0 = v_11542_0 | v_11543_0;
  assign v_11542_0 = v_607_0 ? v_1404_0 : 3'h0;
  assign v_11543_0 = v_26_0 ? v_1390_0 : 3'h0;
  assign v_11544_0 = v_601_0 ? v_1383_0 : 3'h0;
  assign v_11545_0 = v_11546_0 | v_11547_0;
  assign v_11546_0 = v_607_0 ? v_1397_0 : 3'h0;
  assign v_11547_0 = v_26_0 ? v_1383_0 : 3'h0;
  assign v_11548_0 = v_601_0 ? v_1376_0 : 3'h0;
  assign v_11549_0 = v_11550_0 | v_11551_0;
  assign v_11550_0 = v_607_0 ? v_1390_0 : 3'h0;
  assign v_11551_0 = v_26_0 ? v_1376_0 : 3'h0;
  assign v_11552_0 = v_601_0 ? v_1369_0 : 3'h0;
  assign v_11553_0 = v_11554_0 | v_11555_0;
  assign v_11554_0 = v_607_0 ? v_1383_0 : 3'h0;
  assign v_11555_0 = v_26_0 ? v_1369_0 : 3'h0;
  assign v_11556_0 = v_601_0 ? v_1362_0 : 3'h0;
  assign v_11557_0 = v_11558_0 | v_11559_0;
  assign v_11558_0 = v_607_0 ? v_1376_0 : 3'h0;
  assign v_11559_0 = v_26_0 ? v_1362_0 : 3'h0;
  assign v_11560_0 = v_601_0 ? v_1355_0 : 3'h0;
  assign v_11561_0 = v_11562_0 | v_11563_0;
  assign v_11562_0 = v_607_0 ? v_1369_0 : 3'h0;
  assign v_11563_0 = v_26_0 ? v_1355_0 : 3'h0;
  assign v_11564_0 = v_601_0 ? v_1348_0 : 3'h0;
  assign v_11565_0 = v_11566_0 | v_11567_0;
  assign v_11566_0 = v_607_0 ? v_1362_0 : 3'h0;
  assign v_11567_0 = v_26_0 ? v_1348_0 : 3'h0;
  assign v_11568_0 = v_601_0 ? v_1341_0 : 3'h0;
  assign v_11569_0 = v_11570_0 | v_11571_0;
  assign v_11570_0 = v_607_0 ? v_1355_0 : 3'h0;
  assign v_11571_0 = v_26_0 ? v_1341_0 : 3'h0;
  assign v_11572_0 = v_601_0 ? v_1334_0 : 3'h0;
  assign v_11573_0 = v_11574_0 | v_11575_0;
  assign v_11574_0 = v_607_0 ? v_1348_0 : 3'h0;
  assign v_11575_0 = v_26_0 ? v_1334_0 : 3'h0;
  assign v_11576_0 = v_601_0 ? v_1327_0 : 3'h0;
  assign v_11577_0 = v_11578_0 | v_11579_0;
  assign v_11578_0 = v_607_0 ? v_1341_0 : 3'h0;
  assign v_11579_0 = v_26_0 ? v_1327_0 : 3'h0;
  assign v_11580_0 = v_601_0 ? v_1320_0 : 3'h0;
  assign v_11581_0 = v_11582_0 | v_11583_0;
  assign v_11582_0 = v_607_0 ? v_1334_0 : 3'h0;
  assign v_11583_0 = v_26_0 ? v_1320_0 : 3'h0;
  assign v_11584_0 = v_601_0 ? v_1313_0 : 3'h0;
  assign v_11585_0 = v_11586_0 | v_11587_0;
  assign v_11586_0 = v_607_0 ? v_1327_0 : 3'h0;
  assign v_11587_0 = v_26_0 ? v_1313_0 : 3'h0;
  assign v_11588_0 = v_601_0 ? v_1306_0 : 3'h0;
  assign v_11589_0 = v_11590_0 | v_11591_0;
  assign v_11590_0 = v_607_0 ? v_1320_0 : 3'h0;
  assign v_11591_0 = v_26_0 ? v_1306_0 : 3'h0;
  assign v_11592_0 = v_601_0 ? v_1299_0 : 3'h0;
  assign v_11593_0 = v_11594_0 | v_11595_0;
  assign v_11594_0 = v_607_0 ? v_1313_0 : 3'h0;
  assign v_11595_0 = v_26_0 ? v_1299_0 : 3'h0;
  assign v_11596_0 = v_601_0 ? v_1292_0 : 3'h0;
  assign v_11597_0 = v_11598_0 | v_11599_0;
  assign v_11598_0 = v_607_0 ? v_1306_0 : 3'h0;
  assign v_11599_0 = v_26_0 ? v_1292_0 : 3'h0;
  assign v_11600_0 = v_601_0 ? v_1285_0 : 3'h0;
  assign v_11601_0 = v_11602_0 | v_11603_0;
  assign v_11602_0 = v_607_0 ? v_1299_0 : 3'h0;
  assign v_11603_0 = v_26_0 ? v_1285_0 : 3'h0;
  assign v_11604_0 = v_601_0 ? v_1278_0 : 3'h0;
  assign v_11605_0 = v_11606_0 | v_11607_0;
  assign v_11606_0 = v_607_0 ? v_1292_0 : 3'h0;
  assign v_11607_0 = v_26_0 ? v_1278_0 : 3'h0;
  assign v_11608_0 = v_601_0 ? v_1271_0 : 3'h0;
  assign v_11609_0 = v_11610_0 | v_11611_0;
  assign v_11610_0 = v_607_0 ? v_1285_0 : 3'h0;
  assign v_11611_0 = v_26_0 ? v_1271_0 : 3'h0;
  assign v_11612_0 = v_601_0 ? v_1264_0 : 3'h0;
  assign v_11613_0 = v_11614_0 | v_11615_0;
  assign v_11614_0 = v_607_0 ? v_1278_0 : 3'h0;
  assign v_11615_0 = v_26_0 ? v_1264_0 : 3'h0;
  assign v_11616_0 = v_601_0 ? v_1257_0 : 3'h0;
  assign v_11617_0 = v_11618_0 | v_11619_0;
  assign v_11618_0 = v_607_0 ? v_1271_0 : 3'h0;
  assign v_11619_0 = v_26_0 ? v_1257_0 : 3'h0;
  assign v_11620_0 = v_601_0 ? v_1250_0 : 3'h0;
  assign v_11621_0 = v_11622_0 | v_11623_0;
  assign v_11622_0 = v_607_0 ? v_1264_0 : 3'h0;
  assign v_11623_0 = v_26_0 ? v_1250_0 : 3'h0;
  assign v_11624_0 = v_601_0 ? v_1243_0 : 3'h0;
  assign v_11625_0 = v_11626_0 | v_11627_0;
  assign v_11626_0 = v_607_0 ? v_1257_0 : 3'h0;
  assign v_11627_0 = v_26_0 ? v_1243_0 : 3'h0;
  assign v_11628_0 = v_601_0 ? v_1236_0 : 3'h0;
  assign v_11629_0 = v_11630_0 | v_11631_0;
  assign v_11630_0 = v_607_0 ? v_1250_0 : 3'h0;
  assign v_11631_0 = v_26_0 ? v_1236_0 : 3'h0;
  assign v_11632_0 = v_601_0 ? v_1229_0 : 3'h0;
  assign v_11633_0 = v_11634_0 | v_11635_0;
  assign v_11634_0 = v_607_0 ? v_1243_0 : 3'h0;
  assign v_11635_0 = v_26_0 ? v_1229_0 : 3'h0;
  assign v_11636_0 = v_601_0 ? v_1222_0 : 3'h0;
  assign v_11637_0 = v_11638_0 | v_11639_0;
  assign v_11638_0 = v_607_0 ? v_1236_0 : 3'h0;
  assign v_11639_0 = v_26_0 ? v_1222_0 : 3'h0;
  assign v_11640_0 = v_601_0 ? v_1215_0 : 3'h0;
  assign v_11641_0 = v_11642_0 | v_11643_0;
  assign v_11642_0 = v_607_0 ? v_1229_0 : 3'h0;
  assign v_11643_0 = v_26_0 ? v_1215_0 : 3'h0;
  assign v_11644_0 = v_601_0 ? v_1208_0 : 3'h0;
  assign v_11645_0 = v_11646_0 | v_11647_0;
  assign v_11646_0 = v_607_0 ? v_1222_0 : 3'h0;
  assign v_11647_0 = v_26_0 ? v_1208_0 : 3'h0;
  assign v_11648_0 = v_601_0 ? v_1201_0 : 3'h0;
  assign v_11649_0 = v_11650_0 | v_11651_0;
  assign v_11650_0 = v_607_0 ? v_1215_0 : 3'h0;
  assign v_11651_0 = v_26_0 ? v_1201_0 : 3'h0;
  assign v_11652_0 = v_601_0 ? v_1194_0 : 3'h0;
  assign v_11653_0 = v_11654_0 | v_11655_0;
  assign v_11654_0 = v_607_0 ? v_1208_0 : 3'h0;
  assign v_11655_0 = v_26_0 ? v_1194_0 : 3'h0;
  assign v_11656_0 = v_601_0 ? v_1187_0 : 3'h0;
  assign v_11657_0 = v_11658_0 | v_11659_0;
  assign v_11658_0 = v_607_0 ? v_1201_0 : 3'h0;
  assign v_11659_0 = v_26_0 ? v_1187_0 : 3'h0;
  assign v_11660_0 = v_601_0 ? v_1180_0 : 3'h0;
  assign v_11661_0 = v_11662_0 | v_11663_0;
  assign v_11662_0 = v_607_0 ? v_1194_0 : 3'h0;
  assign v_11663_0 = v_26_0 ? v_1180_0 : 3'h0;
  assign v_11664_0 = v_601_0 ? v_1173_0 : 3'h0;
  assign v_11665_0 = v_11666_0 | v_11667_0;
  assign v_11666_0 = v_607_0 ? v_1187_0 : 3'h0;
  assign v_11667_0 = v_26_0 ? v_1173_0 : 3'h0;
  assign v_11668_0 = v_601_0 ? v_1166_0 : 3'h0;
  assign v_11669_0 = v_11670_0 | v_11671_0;
  assign v_11670_0 = v_607_0 ? v_1180_0 : 3'h0;
  assign v_11671_0 = v_26_0 ? v_1166_0 : 3'h0;
  assign v_11672_0 = v_601_0 ? v_1159_0 : 3'h0;
  assign v_11673_0 = v_11674_0 | v_11675_0;
  assign v_11674_0 = v_607_0 ? v_1173_0 : 3'h0;
  assign v_11675_0 = v_26_0 ? v_1159_0 : 3'h0;
  assign v_11676_0 = v_601_0 ? v_1152_0 : 3'h0;
  assign v_11677_0 = v_11678_0 | v_11679_0;
  assign v_11678_0 = v_607_0 ? v_1166_0 : 3'h0;
  assign v_11679_0 = v_26_0 ? v_1152_0 : 3'h0;
  assign v_11680_0 = v_601_0 ? v_1145_0 : 3'h0;
  assign v_11681_0 = v_11682_0 | v_11683_0;
  assign v_11682_0 = v_607_0 ? v_1159_0 : 3'h0;
  assign v_11683_0 = v_26_0 ? v_1145_0 : 3'h0;
  assign v_11684_0 = v_601_0 ? v_1138_0 : 3'h0;
  assign v_11685_0 = v_11686_0 | v_11687_0;
  assign v_11686_0 = v_607_0 ? v_1152_0 : 3'h0;
  assign v_11687_0 = v_26_0 ? v_1138_0 : 3'h0;
  assign v_11688_0 = v_601_0 ? v_1131_0 : 3'h0;
  assign v_11689_0 = v_11690_0 | v_11691_0;
  assign v_11690_0 = v_607_0 ? v_1145_0 : 3'h0;
  assign v_11691_0 = v_26_0 ? v_1131_0 : 3'h0;
  assign v_11692_0 = v_601_0 ? v_1124_0 : 3'h0;
  assign v_11693_0 = v_11694_0 | v_11695_0;
  assign v_11694_0 = v_607_0 ? v_1138_0 : 3'h0;
  assign v_11695_0 = v_26_0 ? v_1124_0 : 3'h0;
  assign v_11696_0 = v_601_0 ? v_1117_0 : 3'h0;
  assign v_11697_0 = v_11698_0 | v_11699_0;
  assign v_11698_0 = v_607_0 ? v_1131_0 : 3'h0;
  assign v_11699_0 = v_26_0 ? v_1117_0 : 3'h0;
  assign v_11700_0 = v_601_0 ? v_1110_0 : 3'h0;
  assign v_11701_0 = v_11702_0 | v_11703_0;
  assign v_11702_0 = v_607_0 ? v_1124_0 : 3'h0;
  assign v_11703_0 = v_26_0 ? v_1110_0 : 3'h0;
  assign v_11704_0 = v_601_0 ? v_1103_0 : 3'h0;
  assign v_11705_0 = v_11706_0 | v_11707_0;
  assign v_11706_0 = v_607_0 ? v_1117_0 : 3'h0;
  assign v_11707_0 = v_26_0 ? v_1103_0 : 3'h0;
  assign v_11708_0 = v_601_0 ? v_1096_0 : 3'h0;
  assign v_11709_0 = v_11710_0 | v_11711_0;
  assign v_11710_0 = v_607_0 ? v_1110_0 : 3'h0;
  assign v_11711_0 = v_26_0 ? v_1096_0 : 3'h0;
  assign v_11712_0 = v_601_0 ? v_1089_0 : 3'h0;
  assign v_11713_0 = v_11714_0 | v_11715_0;
  assign v_11714_0 = v_607_0 ? v_1103_0 : 3'h0;
  assign v_11715_0 = v_26_0 ? v_1089_0 : 3'h0;
  assign v_11716_0 = v_601_0 ? v_1082_0 : 3'h0;
  assign v_11717_0 = v_11718_0 | v_11719_0;
  assign v_11718_0 = v_607_0 ? v_1096_0 : 3'h0;
  assign v_11719_0 = v_26_0 ? v_1082_0 : 3'h0;
  assign v_11720_0 = v_601_0 ? v_1075_0 : 3'h0;
  assign v_11721_0 = v_11722_0 | v_11723_0;
  assign v_11722_0 = v_607_0 ? v_1089_0 : 3'h0;
  assign v_11723_0 = v_26_0 ? v_1075_0 : 3'h0;
  assign v_11724_0 = v_601_0 ? v_1068_0 : 3'h0;
  assign v_11725_0 = v_11726_0 | v_11727_0;
  assign v_11726_0 = v_607_0 ? v_1082_0 : 3'h0;
  assign v_11727_0 = v_26_0 ? v_1068_0 : 3'h0;
  assign v_11728_0 = v_601_0 ? v_1061_0 : 3'h0;
  assign v_11729_0 = v_11730_0 | v_11731_0;
  assign v_11730_0 = v_607_0 ? v_1075_0 : 3'h0;
  assign v_11731_0 = v_26_0 ? v_1061_0 : 3'h0;
  assign v_11732_0 = v_601_0 ? v_1054_0 : 3'h0;
  assign v_11733_0 = v_11734_0 | v_11735_0;
  assign v_11734_0 = v_607_0 ? v_1068_0 : 3'h0;
  assign v_11735_0 = v_26_0 ? v_1054_0 : 3'h0;
  assign v_11736_0 = v_601_0 ? v_1047_0 : 3'h0;
  assign v_11737_0 = v_11738_0 | v_11739_0;
  assign v_11738_0 = v_607_0 ? v_1061_0 : 3'h0;
  assign v_11739_0 = v_26_0 ? v_1047_0 : 3'h0;
  assign v_11740_0 = v_601_0 ? v_1040_0 : 3'h0;
  assign v_11741_0 = v_11742_0 | v_11743_0;
  assign v_11742_0 = v_607_0 ? v_1054_0 : 3'h0;
  assign v_11743_0 = v_26_0 ? v_1040_0 : 3'h0;
  assign v_11744_0 = v_601_0 ? v_1033_0 : 3'h0;
  assign v_11745_0 = v_11746_0 | v_11747_0;
  assign v_11746_0 = v_607_0 ? v_1047_0 : 3'h0;
  assign v_11747_0 = v_26_0 ? v_1033_0 : 3'h0;
  assign v_11748_0 = v_601_0 ? v_1026_0 : 3'h0;
  assign v_11749_0 = v_11750_0 | v_11751_0;
  assign v_11750_0 = v_607_0 ? v_1040_0 : 3'h0;
  assign v_11751_0 = v_26_0 ? v_1026_0 : 3'h0;
  assign v_11752_0 = v_601_0 ? v_1019_0 : 3'h0;
  assign v_11753_0 = v_11754_0 | v_11755_0;
  assign v_11754_0 = v_607_0 ? v_1033_0 : 3'h0;
  assign v_11755_0 = v_26_0 ? v_1019_0 : 3'h0;
  assign v_11756_0 = v_601_0 ? v_1012_0 : 3'h0;
  assign v_11757_0 = v_11758_0 | v_11759_0;
  assign v_11758_0 = v_607_0 ? v_1026_0 : 3'h0;
  assign v_11759_0 = v_26_0 ? v_1012_0 : 3'h0;
  assign v_11760_0 = v_601_0 ? v_1005_0 : 3'h0;
  assign v_11761_0 = v_11762_0 | v_11763_0;
  assign v_11762_0 = v_607_0 ? v_1019_0 : 3'h0;
  assign v_11763_0 = v_26_0 ? v_1005_0 : 3'h0;
  assign v_11764_0 = v_601_0 ? v_998_0 : 3'h0;
  assign v_11765_0 = v_11766_0 | v_11767_0;
  assign v_11766_0 = v_607_0 ? v_1012_0 : 3'h0;
  assign v_11767_0 = v_26_0 ? v_998_0 : 3'h0;
  assign v_11768_0 = v_601_0 ? v_991_0 : 3'h0;
  assign v_11769_0 = v_11770_0 | v_11771_0;
  assign v_11770_0 = v_607_0 ? v_1005_0 : 3'h0;
  assign v_11771_0 = v_26_0 ? v_991_0 : 3'h0;
  assign v_11772_0 = v_601_0 ? v_984_0 : 3'h0;
  assign v_11773_0 = v_11774_0 | v_11775_0;
  assign v_11774_0 = v_607_0 ? v_998_0 : 3'h0;
  assign v_11775_0 = v_26_0 ? v_984_0 : 3'h0;
  assign v_11776_0 = v_601_0 ? v_977_0 : 3'h0;
  assign v_11777_0 = v_11778_0 | v_11779_0;
  assign v_11778_0 = v_607_0 ? v_991_0 : 3'h0;
  assign v_11779_0 = v_26_0 ? v_977_0 : 3'h0;
  assign v_11780_0 = v_601_0 ? v_970_0 : 3'h0;
  assign v_11781_0 = v_11782_0 | v_11783_0;
  assign v_11782_0 = v_607_0 ? v_984_0 : 3'h0;
  assign v_11783_0 = v_26_0 ? v_970_0 : 3'h0;
  assign v_11784_0 = v_601_0 ? v_963_0 : 3'h0;
  assign v_11785_0 = v_11786_0 | v_11787_0;
  assign v_11786_0 = v_607_0 ? v_977_0 : 3'h0;
  assign v_11787_0 = v_26_0 ? v_963_0 : 3'h0;
  assign v_11788_0 = v_601_0 ? v_956_0 : 3'h0;
  assign v_11789_0 = v_11790_0 | v_11791_0;
  assign v_11790_0 = v_607_0 ? v_970_0 : 3'h0;
  assign v_11791_0 = v_26_0 ? v_956_0 : 3'h0;
  assign v_11792_0 = v_601_0 ? v_949_0 : 3'h0;
  assign v_11793_0 = v_11794_0 | v_11795_0;
  assign v_11794_0 = v_607_0 ? v_963_0 : 3'h0;
  assign v_11795_0 = v_26_0 ? v_949_0 : 3'h0;
  assign v_11796_0 = v_601_0 ? v_942_0 : 3'h0;
  assign v_11797_0 = v_11798_0 | v_11799_0;
  assign v_11798_0 = v_607_0 ? v_956_0 : 3'h0;
  assign v_11799_0 = v_26_0 ? v_942_0 : 3'h0;
  assign v_11800_0 = v_601_0 ? v_935_0 : 3'h0;
  assign v_11801_0 = v_11802_0 | v_11803_0;
  assign v_11802_0 = v_607_0 ? v_949_0 : 3'h0;
  assign v_11803_0 = v_26_0 ? v_935_0 : 3'h0;
  assign v_11804_0 = v_601_0 ? v_928_0 : 3'h0;
  assign v_11805_0 = v_11806_0 | v_11807_0;
  assign v_11806_0 = v_607_0 ? v_942_0 : 3'h0;
  assign v_11807_0 = v_26_0 ? v_928_0 : 3'h0;
  assign v_11808_0 = v_601_0 ? v_921_0 : 3'h0;
  assign v_11809_0 = v_11810_0 | v_11811_0;
  assign v_11810_0 = v_607_0 ? v_935_0 : 3'h0;
  assign v_11811_0 = v_26_0 ? v_921_0 : 3'h0;
  assign v_11812_0 = v_601_0 ? v_914_0 : 3'h0;
  assign v_11813_0 = v_11814_0 | v_11815_0;
  assign v_11814_0 = v_607_0 ? v_928_0 : 3'h0;
  assign v_11815_0 = v_26_0 ? v_914_0 : 3'h0;
  assign v_11816_0 = v_601_0 ? v_907_0 : 3'h0;
  assign v_11817_0 = v_11818_0 | v_11819_0;
  assign v_11818_0 = v_607_0 ? v_921_0 : 3'h0;
  assign v_11819_0 = v_26_0 ? v_907_0 : 3'h0;
  assign v_11820_0 = v_601_0 ? v_900_0 : 3'h0;
  assign v_11821_0 = v_11822_0 | v_11823_0;
  assign v_11822_0 = v_607_0 ? v_914_0 : 3'h0;
  assign v_11823_0 = v_26_0 ? v_900_0 : 3'h0;
  assign v_11824_0 = v_601_0 ? v_893_0 : 3'h0;
  assign v_11825_0 = v_11826_0 | v_11827_0;
  assign v_11826_0 = v_607_0 ? v_907_0 : 3'h0;
  assign v_11827_0 = v_26_0 ? v_893_0 : 3'h0;
  assign v_11828_0 = v_601_0 ? v_886_0 : 3'h0;
  assign v_11829_0 = v_11830_0 | v_11831_0;
  assign v_11830_0 = v_607_0 ? v_900_0 : 3'h0;
  assign v_11831_0 = v_26_0 ? v_886_0 : 3'h0;
  assign v_11832_0 = v_601_0 ? v_879_0 : 3'h0;
  assign v_11833_0 = v_11834_0 | v_11835_0;
  assign v_11834_0 = v_607_0 ? v_893_0 : 3'h0;
  assign v_11835_0 = v_26_0 ? v_879_0 : 3'h0;
  assign v_11836_0 = v_601_0 ? v_872_0 : 3'h0;
  assign v_11837_0 = v_11838_0 | v_11839_0;
  assign v_11838_0 = v_607_0 ? v_886_0 : 3'h0;
  assign v_11839_0 = v_26_0 ? v_872_0 : 3'h0;
  assign v_11840_0 = v_601_0 ? v_865_0 : 3'h0;
  assign v_11841_0 = v_11842_0 | v_11843_0;
  assign v_11842_0 = v_607_0 ? v_879_0 : 3'h0;
  assign v_11843_0 = v_26_0 ? v_865_0 : 3'h0;
  assign v_11844_0 = v_601_0 ? v_858_0 : 3'h0;
  assign v_11845_0 = v_11846_0 | v_11847_0;
  assign v_11846_0 = v_607_0 ? v_872_0 : 3'h0;
  assign v_11847_0 = v_26_0 ? v_858_0 : 3'h0;
  assign v_11848_0 = v_601_0 ? v_851_0 : 3'h0;
  assign v_11849_0 = v_11850_0 | v_11851_0;
  assign v_11850_0 = v_607_0 ? v_865_0 : 3'h0;
  assign v_11851_0 = v_26_0 ? v_851_0 : 3'h0;
  assign v_11852_0 = v_601_0 ? v_844_0 : 3'h0;
  assign v_11853_0 = v_11854_0 | v_11855_0;
  assign v_11854_0 = v_607_0 ? v_858_0 : 3'h0;
  assign v_11855_0 = v_26_0 ? v_844_0 : 3'h0;
  assign v_11856_0 = v_601_0 ? v_837_0 : 3'h0;
  assign v_11857_0 = v_11858_0 | v_11859_0;
  assign v_11858_0 = v_607_0 ? v_851_0 : 3'h0;
  assign v_11859_0 = v_26_0 ? v_837_0 : 3'h0;
  assign v_11860_0 = v_601_0 ? v_830_0 : 3'h0;
  assign v_11861_0 = v_11862_0 | v_11863_0;
  assign v_11862_0 = v_607_0 ? v_844_0 : 3'h0;
  assign v_11863_0 = v_26_0 ? v_830_0 : 3'h0;
  assign v_11864_0 = v_601_0 ? v_823_0 : 3'h0;
  assign v_11865_0 = v_11866_0 | v_11867_0;
  assign v_11866_0 = v_607_0 ? v_837_0 : 3'h0;
  assign v_11867_0 = v_26_0 ? v_823_0 : 3'h0;
  assign v_11868_0 = v_601_0 ? v_816_0 : 3'h0;
  assign v_11869_0 = v_11870_0 | v_11871_0;
  assign v_11870_0 = v_607_0 ? v_830_0 : 3'h0;
  assign v_11871_0 = v_26_0 ? v_816_0 : 3'h0;
  assign v_11872_0 = v_601_0 ? v_809_0 : 3'h0;
  assign v_11873_0 = v_11874_0 | v_11875_0;
  assign v_11874_0 = v_607_0 ? v_823_0 : 3'h0;
  assign v_11875_0 = v_26_0 ? v_809_0 : 3'h0;
  assign v_11876_0 = v_601_0 ? v_802_0 : 3'h0;
  assign v_11877_0 = v_11878_0 | v_11879_0;
  assign v_11878_0 = v_607_0 ? v_816_0 : 3'h0;
  assign v_11879_0 = v_26_0 ? v_802_0 : 3'h0;
  assign v_11880_0 = v_601_0 ? v_795_0 : 3'h0;
  assign v_11881_0 = v_11882_0 | v_11883_0;
  assign v_11882_0 = v_607_0 ? v_809_0 : 3'h0;
  assign v_11883_0 = v_26_0 ? v_795_0 : 3'h0;
  assign v_11884_0 = v_601_0 ? v_788_0 : 3'h0;
  assign v_11885_0 = v_11886_0 | v_11887_0;
  assign v_11886_0 = v_607_0 ? v_802_0 : 3'h0;
  assign v_11887_0 = v_26_0 ? v_788_0 : 3'h0;
  assign v_11888_0 = v_601_0 ? v_781_0 : 3'h0;
  assign v_11889_0 = v_11890_0 | v_11891_0;
  assign v_11890_0 = v_607_0 ? v_795_0 : 3'h0;
  assign v_11891_0 = v_26_0 ? v_781_0 : 3'h0;
  assign v_11892_0 = v_601_0 ? v_774_0 : 3'h0;
  assign v_11893_0 = v_11894_0 | v_11895_0;
  assign v_11894_0 = v_607_0 ? v_788_0 : 3'h0;
  assign v_11895_0 = v_26_0 ? v_774_0 : 3'h0;
  assign v_11896_0 = v_601_0 ? v_767_0 : 3'h0;
  assign v_11897_0 = v_11898_0 | v_11899_0;
  assign v_11898_0 = v_607_0 ? v_781_0 : 3'h0;
  assign v_11899_0 = v_26_0 ? v_767_0 : 3'h0;
  assign v_11900_0 = v_601_0 ? v_760_0 : 3'h0;
  assign v_11901_0 = v_11902_0 | v_11903_0;
  assign v_11902_0 = v_607_0 ? v_774_0 : 3'h0;
  assign v_11903_0 = v_26_0 ? v_760_0 : 3'h0;
  assign v_11904_0 = v_601_0 ? v_753_0 : 3'h0;
  assign v_11905_0 = v_11906_0 | v_11907_0;
  assign v_11906_0 = v_607_0 ? v_767_0 : 3'h0;
  assign v_11907_0 = v_26_0 ? v_753_0 : 3'h0;
  assign v_11908_0 = v_601_0 ? v_746_0 : 3'h0;
  assign v_11909_0 = v_11910_0 | v_11911_0;
  assign v_11910_0 = v_607_0 ? v_760_0 : 3'h0;
  assign v_11911_0 = v_26_0 ? v_746_0 : 3'h0;
  assign v_11912_0 = v_601_0 ? v_739_0 : 3'h0;
  assign v_11913_0 = v_11914_0 | v_11915_0;
  assign v_11914_0 = v_607_0 ? v_753_0 : 3'h0;
  assign v_11915_0 = v_26_0 ? v_739_0 : 3'h0;
  assign v_11916_0 = v_601_0 ? v_732_0 : 3'h0;
  assign v_11917_0 = v_11918_0 | v_11919_0;
  assign v_11918_0 = v_607_0 ? v_746_0 : 3'h0;
  assign v_11919_0 = v_26_0 ? v_732_0 : 3'h0;
  assign v_11920_0 = v_601_0 ? v_725_0 : 3'h0;
  assign v_11921_0 = v_11922_0 | v_11923_0;
  assign v_11922_0 = v_607_0 ? v_739_0 : 3'h0;
  assign v_11923_0 = v_26_0 ? v_725_0 : 3'h0;
  assign v_11924_0 = v_601_0 ? v_718_0 : 3'h0;
  assign v_11925_0 = v_11926_0 | v_11927_0;
  assign v_11926_0 = v_607_0 ? v_732_0 : 3'h0;
  assign v_11927_0 = v_26_0 ? v_718_0 : 3'h0;
  assign v_11928_0 = v_601_0 ? v_711_0 : 3'h0;
  assign v_11929_0 = v_11930_0 | v_11931_0;
  assign v_11930_0 = v_607_0 ? v_725_0 : 3'h0;
  assign v_11931_0 = v_26_0 ? v_711_0 : 3'h0;
  assign v_11932_0 = v_601_0 ? v_704_0 : 3'h0;
  assign v_11933_0 = v_11934_0 | v_11935_0;
  assign v_11934_0 = v_607_0 ? v_718_0 : 3'h0;
  assign v_11935_0 = v_26_0 ? v_704_0 : 3'h0;
  assign v_11936_0 = v_601_0 ? v_697_0 : 3'h0;
  assign v_11937_0 = v_11938_0 | v_11939_0;
  assign v_11938_0 = v_607_0 ? v_711_0 : 3'h0;
  assign v_11939_0 = v_26_0 ? v_697_0 : 3'h0;
  assign v_11940_0 = v_601_0 ? v_690_0 : 3'h0;
  assign v_11941_0 = v_11942_0 | v_11943_0;
  assign v_11942_0 = v_607_0 ? v_704_0 : 3'h0;
  assign v_11943_0 = v_26_0 ? v_690_0 : 3'h0;
  assign v_11944_0 = v_601_0 ? v_50_0 : 3'h0;
  assign v_11945_0 = v_11946_0 | v_11947_0;
  assign v_11946_0 = v_607_0 ? v_697_0 : 3'h0;
  assign v_11947_0 = v_26_0 ? v_50_0 : 3'h0;
  assign v_11949_0 = v_11950_0 | v_11951_0;
  assign v_11950_0 = v_614_0 | v_656_0;
  assign v_11951_0 = v_11952_0 | v_11953_0;
  assign v_11952_0 = v_589_0 | v_601_0;
  assign v_11953_0 = v_607_0 | v_26_0;
  assign v_11954_0 = v_11955_0 | v_12053_0;
  assign v_11955_0 = v_11956_0 | v_12052_0;
  assign v_11956_0 = v_614_0 ? v_11957_0 : 3'h0;
  assign v_11957_0 = v_11958_0 ? v_12002_0 : v_12013_0;
  assign v_11958_0 = v_11959_0 & v_11964_0;
  assign v_11959_0 = v_11960_0 & v_11961_0;
  assign _act_11962_0 = v_656_0 | v_11963_0;
  assign v_11963_0 = v_601_0 | v_26_0;
  assign v_11964_0 = v_11965_0 == v_11993_0;
  assign v_11966_0 = v_11967_0 | v_11991_0;
  assign v_11967_0 = 1'h1 ? v_11968_0 : 10'h0;
  assign v_11968_0 = _act_11969_0 ? v_11974_0 : v_11989_0;
  assign _act_11969_0 = v_11970_0 | v_11971_0;
  assign v_11970_0 = v_614_0 | v_656_0;
  assign v_11971_0 = v_11972_0 | v_11973_0;
  assign v_11972_0 = v_589_0 | v_601_0;
  assign v_11973_0 = v_607_0 | v_26_0;
  assign v_11974_0 = v_11975_0 | v_11982_0;
  assign v_11975_0 = v_11976_0 | v_11978_0;
  assign v_11976_0 = v_11977_0 ? v_597_0 : 10'h0;
  assign v_11977_0 = ~_act_11969_0;
  assign v_11978_0 = v_11979_0 | v_11981_0;
  assign v_11979_0 = v_589_0 ? v_11980_0 : 10'h0;
  assign v_11980_0 = v_597_0 - 10'h1;
  assign v_11981_0 = v_601_0 ? v_597_0 : 10'h0;
  assign v_11982_0 = v_11983_0 | v_11986_0;
  assign v_11983_0 = v_11984_0 | v_11985_0;
  assign v_11984_0 = v_607_0 ? v_11980_0 : 10'h0;
  assign v_11985_0 = v_26_0 ? v_597_0 : 10'h0;
  assign v_11986_0 = v_11987_0 | v_11988_0;
  assign v_11987_0 = v_614_0 ? v_11980_0 : 10'h0;
  assign v_11988_0 = v_656_0 ? v_597_0 : 10'h0;
  assign v_11990_0 = _act_11969_0 & 1'h1;
  assign v_11991_0 = v_11992_0 ? 10'bxxxxxxxxxx : 10'h0;
  assign v_11992_0 = ~1'h1;
  assign v_11994_0 = v_11995_0 | v_11998_0;
  assign v_11995_0 = v_11996_0 | v_11997_0;
  assign v_11996_0 = v_601_0 ? v_597_0 : 10'h0;
  assign v_11997_0 = v_26_0 ? v_597_0 : 10'h0;
  assign v_11998_0 = v_11999_0 | v_12000_0;
  assign v_11999_0 = v_656_0 ? v_597_0 : 10'h0;
  assign v_12000_0 = v_12001_0 ? 10'bxxxxxxxxxx : 10'h0;
  assign v_12001_0 = ~_act_11962_0;
  assign v_12003_0 = v_12004_0 | v_12007_0;
  assign v_12004_0 = v_12005_0 | v_12006_0;
  assign v_12005_0 = v_601_0 ? v_11948_0 : 3'h0;
  assign v_12006_0 = v_26_0 ? v_11948_0 : 3'h0;
  assign v_12007_0 = v_12008_0 | v_12009_0;
  assign v_12008_0 = v_656_0 ? v_11948_0 : 3'h0;
  assign v_12009_0 = v_12010_0 ? 3'bxxx : 3'h0;
  assign v_12010_0 = ~v_12011_0;
  assign v_12011_0 = v_656_0 | v_12012_0;
  assign v_12012_0 = v_601_0 | v_26_0;
  BlockRAMTrueDual#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(3))
    ram12013
      (.CLK(clock),
       .DI_A(v_12018_0),
       .ADDR_A(v_12014_0),
       .WE_A(v_12020_0),
       .DO_A(v_12013_0),
       .DI_B(v_12032_0),
       .ADDR_B(v_12022_0),
       .WE_B(v_12042_0),
       .DO_B(v_12013_1));
  assign v_12014_0 = v_12015_0 | v_12016_0;
  assign v_12015_0 = 1'h1 ? v_11968_0 : 10'h0;
  assign v_12016_0 = v_12017_0 ? 10'bxxxxxxxxxx : 10'h0;
  assign v_12017_0 = ~1'h1;
  assign v_12018_0 = v_12019_0 ? 3'bxxx : 3'h0;
  assign v_12019_0 = ~1'h0;
  assign v_12020_0 = v_12021_0 ? 1'h0 : 1'h0;
  assign v_12021_0 = ~1'h0;
  assign v_12022_0 = v_12023_0 | v_12026_0;
  assign v_12023_0 = v_12024_0 | v_12025_0;
  assign v_12024_0 = v_601_0 ? v_597_0 : 10'h0;
  assign v_12025_0 = v_26_0 ? v_597_0 : 10'h0;
  assign v_12026_0 = v_12027_0 | v_12028_0;
  assign v_12027_0 = v_656_0 ? v_597_0 : 10'h0;
  assign v_12028_0 = v_12029_0 ? 10'bxxxxxxxxxx : 10'h0;
  assign v_12029_0 = ~v_12030_0;
  assign v_12030_0 = v_656_0 | v_12031_0;
  assign v_12031_0 = v_601_0 | v_26_0;
  assign v_12032_0 = v_12033_0 | v_12036_0;
  assign v_12033_0 = v_12034_0 | v_12035_0;
  assign v_12034_0 = v_601_0 ? v_11948_0 : 3'h0;
  assign v_12035_0 = v_26_0 ? v_11948_0 : 3'h0;
  assign v_12036_0 = v_12037_0 | v_12038_0;
  assign v_12037_0 = v_656_0 ? v_11948_0 : 3'h0;
  assign v_12038_0 = v_12039_0 ? 3'bxxx : 3'h0;
  assign v_12039_0 = ~v_12040_0;
  assign v_12040_0 = v_656_0 | v_12041_0;
  assign v_12041_0 = v_601_0 | v_26_0;
  assign v_12042_0 = v_12043_0 | v_12046_0;
  assign v_12043_0 = v_12044_0 | v_12045_0;
  assign v_12044_0 = v_601_0 ? 1'h1 : 1'h0;
  assign v_12045_0 = v_26_0 ? 1'h1 : 1'h0;
  assign v_12046_0 = v_12047_0 | v_12048_0;
  assign v_12047_0 = v_656_0 ? 1'h1 : 1'h0;
  assign v_12048_0 = v_12049_0 ? 1'h0 : 1'h0;
  assign v_12049_0 = ~v_12050_0;
  assign v_12050_0 = v_656_0 | v_12051_0;
  assign v_12051_0 = v_601_0 | v_26_0;
  assign v_12052_0 = v_656_0 ? v_328_0 : 3'h0;
  assign v_12053_0 = v_12054_0 | v_12057_0;
  assign v_12054_0 = v_12055_0 | v_12056_0;
  assign v_12055_0 = v_589_0 ? v_11957_0 : 3'h0;
  assign v_12056_0 = v_601_0 ? v_50_0 : 3'h0;
  assign v_12057_0 = v_12058_0 | v_12059_0;
  assign v_12058_0 = v_607_0 ? v_11957_0 : 3'h0;
  assign v_12059_0 = v_26_0 ? v_50_0 : 3'h0;
  assign v_12060_0 = v_16_0 & v_12061_0;
  assign v_12061_0 = ~v_12062_0;
  assign v_12062_0 = v_12063_0 | v_12078_0;
  assign v_12063_0 = ~v_12064_0;
  assign v_12064_0 = v_12065_0 & v_7_0;
  assign v_12066_0 = v_12067_0 | v_12069_0;
  assign v_12067_0 = v_12068_0 & v_606_0;
  assign v_12068_0 = v_578_0 == 16'h0;
  assign v_12069_0 = v_12070_0 | v_86_0;
  assign v_12070_0 = v_12071_0 & v_148_0;
  assign v_12071_0 = v_12072_0 & v_94_0;
  assign v_12072_0 = v_578_0 <= v_97_0;
  assign v_12073_0 = v_12074_0 | v_12075_0;
  assign v_12074_0 = v_12067_0 ? 1'h1 : 1'h0;
  assign v_12075_0 = v_12076_0 | v_12077_0;
  assign v_12076_0 = v_12070_0 ? 1'h1 : 1'h0;
  assign v_12077_0 = v_86_0 ? 1'h0 : 1'h0;
  assign v_12079_0 = v_12060_0 | v_88_0;
  assign v_12080_0 = v_12081_0 | v_12082_0;
  assign v_12081_0 = v_12060_0 ? 1'h1 : 1'h0;
  assign v_12082_0 = v_88_0 ? 1'h0 : 1'h0;
  assign v_12083_0 = ~v_12084_0;
  assign v_12084_0 = 16'h5 <= v_12_0;
  assign v_12085_0 = v_12_0 + 16'h1;
  assign v_12087_0 = 1'h1 & v_12088_0;
  assign v_12088_0 = v_12089_0 | v_12146_0;
  assign v_12089_0 = ~v_12090_0;
  assign v_12091_0 = v_12092_0 | _act_12095_0;
  assign v_12093_0 = v_12094_0 | v_12142_0;
  assign v_12094_0 = _act_12095_0 & v_12140_0;
  assign _act_12095_0 = v_12096_0 & 1'h1;
  assign v_12096_0 = v_12097_0 & v_12098_0;
  assign v_12097_0 = ~v_12092_0;
  assign v_12098_0 = ~v_12099_0;
  assign v_12100_0 = v_12101_0 | v_12135_0;
  assign v_12101_0 = v_12102_0 & v_12132_0;
  assign v_12102_0 = v_12103_0 == v_12110_0;
  assign v_12103_0 = v_12104_0 ? v_12108_0 : v_12109_0;
  assign v_12104_0 = v_12105_0 | v_12106_0;
  assign v_12105_0 = _act_12095_0 ? 1'h1 : 1'h0;
  assign v_12106_0 = v_12107_0 ? 1'h0 : 1'h0;
  assign v_12107_0 = ~_act_12095_0;
  assign v_12108_0 = v_12109_0 + 5'h1;
  assign _act_12111_0 = 1'h1 & _act_12112_0;
  assign _act_12112_0 = v_12113_0 | v_12116_0;
  assign v_12113_0 = v_12114_0 | v_12115_0;
  assign v_12114_0 = v_13_0 & v_11_0;
  assign v_12115_0 = v_6_0 & v_11_0;
  assign v_12116_0 = v_12117_0 | v_12126_0;
  assign v_12117_0 = v_12118_0 | v_12119_0;
  assign v_12118_0 = v_147_0 & v_11_0;
  assign v_12119_0 = v_12120_0 & v_11_0;
  assign v_12120_0 = v_12121_0 & v_12124_0;
  assign v_12121_0 = v_86_0 & v_12122_0;
  assign v_12122_0 = ~v_12123_0;
  assign v_12123_0 = v_40_0 & v_45_0;
  assign v_12124_0 = ~v_12125_0;
  assign v_12125_0 = v_40_0 & v_46_0;
  assign v_12126_0 = v_12127_0 | v_12129_0;
  assign v_12127_0 = v_12128_0 & v_11_0;
  assign v_12128_0 = v_12121_0 & v_12125_0;
  assign v_12129_0 = v_12130_0 & v_11_0;
  assign v_12130_0 = v_86_0 & v_12123_0;
  assign v_12131_0 = v_12110_0 + 5'h1;
  assign v_12132_0 = v_12104_0 & v_12133_0;
  assign v_12133_0 = 1'h1 & v_12134_0;
  assign v_12134_0 = ~_act_12112_0;
  assign v_12135_0 = v_12136_0 & _act_12111_0;
  assign v_12136_0 = ~v_12104_0;
  assign v_12137_0 = v_12138_0 | v_12139_0;
  assign v_12138_0 = v_12101_0 ? 1'h1 : 1'h0;
  assign v_12139_0 = v_12135_0 ? 1'h0 : 1'h0;
  assign v_12140_0 = 1'h1 & v_12141_0;
  assign v_12141_0 = ~v_12088_0;
  assign v_12142_0 = v_12092_0 & v_12087_0;
  assign v_12143_0 = v_12144_0 | v_12145_0;
  assign v_12144_0 = v_12094_0 ? 1'h1 : 1'h0;
  assign v_12145_0 = v_12142_0 ? _act_12095_0 : 1'h0;
  assign v_12146_0 = v_12147_0 | v_12152_0;
  assign v_12147_0 = v_12148_0 ? 1'h0 : 1'h0;
  assign v_12148_0 = ~v_12149_0;
  assign v_12149_0 = v_12150_0 | v_12151_0;
  assign v_12150_0 = v_11_0 & v_93_0;
  assign v_12151_0 = v_11_0 & v_6_0;
  assign v_12152_0 = v_12153_0 | v_12154_0;
  assign v_12153_0 = v_12150_0 ? 1'h1 : 1'h0;
  assign v_12154_0 = v_12151_0 ? 1'h1 : 1'h0;
  assign v_12155_0 = v_12092_0 ? v_12156_0 : v_12165_0;
  assign v_12157_0 = v_12158_0 & 1'h1;
  assign v_12158_0 = v_12159_0 | v_12162_0;
  assign v_12159_0 = v_12160_0 ? 1'h0 : 1'h0;
  assign v_12160_0 = ~v_12161_0;
  assign v_12161_0 = v_12094_0 | v_12142_0;
  assign v_12162_0 = v_12163_0 | v_12164_0;
  assign v_12163_0 = v_12094_0 ? 1'h1 : 1'h0;
  assign v_12164_0 = v_12142_0 ? 1'h1 : 1'h0;
  assign v_12165_0 = v_12166_0 | v_12224_0;
  assign v_12166_0 = _act_12095_0 ? v_12167_0 : 16'h0;
  assign v_12167_0 = v_12168_0 ? v_12183_0 : v_12203_0;
  assign v_12168_0 = v_12169_0 & v_12172_0;
  assign v_12169_0 = v_12170_0 & v_12171_0;
  assign v_12172_0 = v_12173_0 == v_12178_0;
  assign v_12174_0 = v_12175_0 | v_12176_0;
  assign v_12175_0 = 1'h1 ? v_12103_0 : 5'h0;
  assign v_12176_0 = v_12177_0 ? 5'bxxxxx : 5'h0;
  assign v_12177_0 = ~1'h1;
  assign v_12179_0 = v_12180_0 | v_12181_0;
  assign v_12180_0 = _act_12111_0 ? v_12110_0 : 5'h0;
  assign v_12181_0 = v_12182_0 ? 5'bxxxxx : 5'h0;
  assign v_12182_0 = ~_act_12111_0;
  assign v_12184_0 = v_12185_0 | v_12201_0;
  assign v_12185_0 = _act_12111_0 ? v_12186_0 : 16'h0;
  assign v_12186_0 = v_12187_0 | v_12193_0;
  assign v_12187_0 = v_12188_0 | v_12190_0;
  assign v_12188_0 = v_12189_0 ? 16'bxxxxxxxxxxxxxxxx : 16'h0;
  assign v_12189_0 = ~_act_12112_0;
  assign v_12190_0 = v_12191_0 | v_12192_0;
  assign v_12191_0 = v_12118_0 ? v_10_0 : 16'h0;
  assign v_12192_0 = v_12119_0 ? v_10_0 : 16'h0;
  assign v_12193_0 = v_12194_0 | v_12198_0;
  assign v_12194_0 = v_12195_0 | v_12197_0;
  assign v_12195_0 = v_12127_0 ? v_12196_0 : 16'h0;
  assign v_12196_0 = v_10_0 + 16'h1;
  assign v_12197_0 = v_12129_0 ? 16'h0 : 16'h0;
  assign v_12198_0 = v_12199_0 | v_12200_0;
  assign v_12199_0 = v_12114_0 ? 16'h0 : 16'h0;
  assign v_12200_0 = v_12115_0 ? v_10_0 : 16'h0;
  assign v_12201_0 = v_12202_0 ? 16'bxxxxxxxxxxxxxxxx : 16'h0;
  assign v_12202_0 = ~_act_12111_0;
  BlockRAMTrueDual#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(5), .DATA_WIDTH(16))
    ram12203
      (.CLK(clock),
       .DI_A(v_12208_0),
       .ADDR_A(v_12204_0),
       .WE_A(v_12210_0),
       .DO_A(v_12203_0),
       .DI_B(v_12216_0),
       .ADDR_B(v_12212_0),
       .WE_B(v_12220_0),
       .DO_B(v_12203_1));
  assign v_12204_0 = v_12205_0 | v_12206_0;
  assign v_12205_0 = 1'h1 ? v_12103_0 : 5'h0;
  assign v_12206_0 = v_12207_0 ? 5'bxxxxx : 5'h0;
  assign v_12207_0 = ~1'h1;
  assign v_12208_0 = v_12209_0 ? 16'bxxxxxxxxxxxxxxxx : 16'h0;
  assign v_12209_0 = ~1'h0;
  assign v_12210_0 = v_12211_0 ? 1'h0 : 1'h0;
  assign v_12211_0 = ~1'h0;
  assign v_12212_0 = v_12213_0 | v_12214_0;
  assign v_12213_0 = _act_12111_0 ? v_12110_0 : 5'h0;
  assign v_12214_0 = v_12215_0 ? 5'bxxxxx : 5'h0;
  assign v_12215_0 = ~_act_12111_0;
  assign v_12216_0 = v_12217_0 | v_12218_0;
  assign v_12217_0 = _act_12111_0 ? v_12186_0 : 16'h0;
  assign v_12218_0 = v_12219_0 ? 16'bxxxxxxxxxxxxxxxx : 16'h0;
  assign v_12219_0 = ~_act_12111_0;
  assign v_12220_0 = v_12221_0 | v_12222_0;
  assign v_12221_0 = _act_12111_0 ? 1'h1 : 1'h0;
  assign v_12222_0 = v_12223_0 ? 1'h0 : 1'h0;
  assign v_12223_0 = ~_act_12111_0;
  assign v_12224_0 = v_12225_0 ? 16'bxxxxxxxxxxxxxxxx : 16'h0;
  assign v_12225_0 = ~_act_12095_0;
  assign v_12227_0 = v_12228_0 | v_12233_0;
  assign v_12228_0 = v_12229_0 | v_12231_0;
  assign v_12229_0 = v_13_0 & v_12230_0;
  assign v_12230_0 = ~v_11_0;
  assign v_12231_0 = v_6_0 & v_12232_0;
  assign v_12232_0 = ~v_11_0;
  assign v_12233_0 = v_12234_0 | v_12239_0;
  assign v_12234_0 = v_12235_0 | v_12237_0;
  assign v_12235_0 = v_147_0 & v_12236_0;
  assign v_12236_0 = ~v_11_0;
  assign v_12237_0 = v_12120_0 & v_12238_0;
  assign v_12238_0 = ~v_11_0;
  assign v_12239_0 = v_12240_0 | v_12242_0;
  assign v_12240_0 = v_12128_0 & v_12241_0;
  assign v_12241_0 = ~v_11_0;
  assign v_12242_0 = v_12130_0 & v_12243_0;
  assign v_12243_0 = ~v_11_0;
  assign v_12244_0 = v_12245_0 | v_12248_0;
  assign v_12245_0 = v_12246_0 | v_12247_0;
  assign v_12246_0 = v_12229_0 ? 16'h0 : 16'h0;
  assign v_12247_0 = v_12231_0 ? v_10_0 : 16'h0;
  assign v_12248_0 = v_12249_0 | v_12252_0;
  assign v_12249_0 = v_12250_0 | v_12251_0;
  assign v_12250_0 = v_12235_0 ? v_10_0 : 16'h0;
  assign v_12251_0 = v_12237_0 ? v_10_0 : 16'h0;
  assign v_12252_0 = v_12253_0 | v_12254_0;
  assign v_12253_0 = v_12240_0 ? v_12196_0 : 16'h0;
  assign v_12254_0 = v_12242_0 ? 16'h0 : 16'h0;
  assign v_12255_0 = v_12256_0 | v_12258_0;
  assign v_12256_0 = 1'h1 & v_12257_0;
  assign v_12257_0 = v_10_0 == 16'h1;
  assign v_12258_0 = v_12259_0 | 1'h0;
  assign v_12259_0 = v_12260_0 & v_12264_0;
  assign v_12260_0 = v_642_0 | v_12261_0;
  assign v_12261_0 = v_12262_0 & v_12263_0;
  assign v_12262_0 = ~v_620_0;
  assign v_12263_0 = ~v_628_0;
  assign v_12264_0 = v_10_0 == 16'h2;
  assign v_12265_0 = ~v_3_0;
  assign v_12266_0 = v_10_0 == 16'h0;
  assign v_12268_0 = v_2_0 & v_6_0;
  assign v_12270_0 = v_2_0 & v_6_0;
  assign v_12272_0 = v_12273_0 & v_6_0;
  assign v_12273_0 = v_3_0 & v_12274_0;
  assign v_12274_0 = v_10_0 == 16'h1;
  assign v_12276_0 = v_12273_0 & v_6_0;
  assign v_12278_0 = v_12279_0 & v_6_0;
  assign v_12279_0 = v_3_0 & v_12280_0;
  assign v_12280_0 = v_10_0 == 16'h2;
  assign v_12282_0 = v_12279_0 & v_6_0;
  assign v_12284_0 = v_12279_0 & v_6_0;
  assign v_12286_0 = v_12287_0 & v_30_0;
  assign v_12287_0 = ~v_12288_0;
  assign v_12289_0 = v_12290_0 ? v_97_0 : v_12_0;
  assign v_12290_0 = v_97_0 != 16'h0;
  assign v_12292_0 = v_34_0 & v_32_0;
  assign v_12295_0 = v_12294_0 + 32'h1;
  assign v_12297_0 = v_14_0 & v_12084_0;
  assign v_12299_0 = v_12300_0 & v_147_0;
  assign v_12300_0 = 1'h0 & v_12301_0;
  assign v_12301_0 = v_10_0 == 16'h0;
  assign v_12303_0 = v_12300_0 & v_147_0;
  assign v_12305_0 = v_12300_0 & v_147_0;
  assign v_12307_0 = v_12308_0 & v_147_0;
  assign v_12308_0 = 1'h0 & v_12309_0;
  assign v_12309_0 = v_10_0 == 16'h1;
  assign v_12311_0 = v_12308_0 & v_147_0;
  assign v_12313_0 = v_12314_0 & v_147_0;
  assign v_12314_0 = 1'h0 & v_12315_0;
  assign v_12315_0 = v_10_0 == 16'h2;
  assign v_12317_0 = v_12314_0 & v_147_0;
  assign v_12319_0 = v_12314_0 & v_147_0;
  assign v_12322_0 = v_20_0 & v_19_0;
  assign v_12324_0 = v_12325_0 & v_19_0;
  assign v_12325_0 = ~v_21_0;
  assign in_consume_en = v_12327_0;
  assign v_12327_0 = v_12328_0 | v_12331_0;
  assign v_12328_0 = v_12329_0 ? 1'h1 : 1'h0;
  assign v_12329_0 = v_12330_0 & 1'h1;
  assign v_12330_0 = in_canPeek;
  assign v_12331_0 = v_12332_0 ? 1'h0 : 1'h0;
  assign v_12332_0 = ~v_12329_0;
  assign out_canPeek = v_12334_0;
  assign v_12335_0 = 1'h1 & v_12336_0;
  assign v_12336_0 = v_12337_0 | v_12338_0;
  assign v_12337_0 = ~v_12334_0;
  assign v_12338_0 = v_12339_0 | v_12342_0;
  assign v_12339_0 = v_12340_0 ? 1'h1 : 1'h0;
  assign v_12340_0 = v_12341_0 & 1'h1;
  assign v_12341_0 = out_consume_en;
  assign v_12342_0 = v_12343_0 ? 1'h0 : 1'h0;
  assign v_12343_0 = ~v_12340_0;
  assign v_12344_0 = v_12345_0 | _act_12348_0;
  assign v_12346_0 = v_12347_0 | v_12351_0;
  assign v_12347_0 = _act_12348_0 & v_12349_0;
  assign _act_12348_0 = v_19_0 | v_12297_0;
  assign v_12349_0 = 1'h1 & v_12350_0;
  assign v_12350_0 = ~v_12336_0;
  assign v_12351_0 = v_12345_0 & v_12335_0;
  assign v_12352_0 = v_12353_0 | v_12354_0;
  assign v_12353_0 = v_12347_0 ? 1'h1 : 1'h0;
  assign v_12354_0 = v_12351_0 ? _act_12348_0 : 1'h0;
  assign out_peek = v_12356_0;
  assign v_12357_0 = v_12345_0 ? v_12358_0 : v_12367_0;
  assign v_12359_0 = v_12360_0 & 1'h1;
  assign v_12360_0 = v_12361_0 | v_12364_0;
  assign v_12361_0 = v_12362_0 ? 1'h0 : 1'h0;
  assign v_12362_0 = ~v_12363_0;
  assign v_12363_0 = v_12347_0 | v_12351_0;
  assign v_12364_0 = v_12365_0 | v_12366_0;
  assign v_12365_0 = v_12347_0 ? 1'h1 : 1'h0;
  assign v_12366_0 = v_12351_0 ? 1'h1 : 1'h0;
  assign v_12367_0 = v_12368_0 | v_12370_0;
  assign v_12368_0 = v_12369_0 ? 8'bxxxxxxxx : 8'h0;
  assign v_12369_0 = ~_act_12348_0;
  assign v_12370_0 = v_12371_0 | v_12372_0;
  assign v_12371_0 = v_19_0 ? 8'h46 : 8'h0;
  assign v_12372_0 = v_12297_0 ? 8'h50 : 8'h0;
  assign v_12373_0 = in_peek;
  // Always block
  //////////////////////////////////////////////////////////////////////////////
  always @(posedge clock) begin
    if (reset) begin
      v_3_0 <= 1'h0;
      v_12_0 <= 16'h0;
      v_18_0 <= 1'h0;
      v_23_0 <= 10'h0;
      v_34_0 <= 1'h1;
      v_40_0 <= 1'h1;
      v_52_0 <= 16'h0;
      v_54_0 <= 3'h0;
      v_58_0 <= 1'h0;
      v_60_0 <= 1'h0;
      v_67_0 <= 1'h1;
      v_77_0 <= 5'h0;
      v_78_0 <= 5'h0;
      v_91_0 <= 1'h0;
      v_97_0 <= 16'h0;
      v_191_0 <= 3'h0;
      v_205_0 <= 1'h0;
      v_206_0 <= 1'h0;
      v_208_0 <= 5'h0;
      v_213_0 <= 5'h0;
      v_218_0 <= 3'h0;
      v_271_0 <= 3'h0;
      v_330_0 <= 16'h0;
      v_332_0 <= 3'h0;
      v_336_0 <= 1'h0;
      v_338_0 <= 1'h0;
      v_345_0 <= 1'h1;
      v_355_0 <= 5'h0;
      v_356_0 <= 5'h0;
      v_434_0 <= 3'h0;
      v_448_0 <= 1'h0;
      v_449_0 <= 1'h0;
      v_451_0 <= 5'h0;
      v_456_0 <= 5'h0;
      v_461_0 <= 3'h0;
      v_514_0 <= 3'h0;
      v_578_0 <= 16'h0;
      v_597_0 <= 10'h0;
      v_615_0 <= 1'h0;
      v_616_0 <= 1'h0;
      v_620_0 <= 1'h0;
      v_642_0 <= 1'h0;
      v_690_0 <= 3'h0;
      v_697_0 <= 3'h0;
      v_704_0 <= 3'h0;
      v_711_0 <= 3'h0;
      v_718_0 <= 3'h0;
      v_725_0 <= 3'h0;
      v_732_0 <= 3'h0;
      v_739_0 <= 3'h0;
      v_746_0 <= 3'h0;
      v_753_0 <= 3'h0;
      v_760_0 <= 3'h0;
      v_767_0 <= 3'h0;
      v_774_0 <= 3'h0;
      v_781_0 <= 3'h0;
      v_788_0 <= 3'h0;
      v_795_0 <= 3'h0;
      v_802_0 <= 3'h0;
      v_809_0 <= 3'h0;
      v_816_0 <= 3'h0;
      v_823_0 <= 3'h0;
      v_830_0 <= 3'h0;
      v_837_0 <= 3'h0;
      v_844_0 <= 3'h0;
      v_851_0 <= 3'h0;
      v_858_0 <= 3'h0;
      v_865_0 <= 3'h0;
      v_872_0 <= 3'h0;
      v_879_0 <= 3'h0;
      v_886_0 <= 3'h0;
      v_893_0 <= 3'h0;
      v_900_0 <= 3'h0;
      v_907_0 <= 3'h0;
      v_914_0 <= 3'h0;
      v_921_0 <= 3'h0;
      v_928_0 <= 3'h0;
      v_935_0 <= 3'h0;
      v_942_0 <= 3'h0;
      v_949_0 <= 3'h0;
      v_956_0 <= 3'h0;
      v_963_0 <= 3'h0;
      v_970_0 <= 3'h0;
      v_977_0 <= 3'h0;
      v_984_0 <= 3'h0;
      v_991_0 <= 3'h0;
      v_998_0 <= 3'h0;
      v_1005_0 <= 3'h0;
      v_1012_0 <= 3'h0;
      v_1019_0 <= 3'h0;
      v_1026_0 <= 3'h0;
      v_1033_0 <= 3'h0;
      v_1040_0 <= 3'h0;
      v_1047_0 <= 3'h0;
      v_1054_0 <= 3'h0;
      v_1061_0 <= 3'h0;
      v_1068_0 <= 3'h0;
      v_1075_0 <= 3'h0;
      v_1082_0 <= 3'h0;
      v_1089_0 <= 3'h0;
      v_1096_0 <= 3'h0;
      v_1103_0 <= 3'h0;
      v_1110_0 <= 3'h0;
      v_1117_0 <= 3'h0;
      v_1124_0 <= 3'h0;
      v_1131_0 <= 3'h0;
      v_1138_0 <= 3'h0;
      v_1145_0 <= 3'h0;
      v_1152_0 <= 3'h0;
      v_1159_0 <= 3'h0;
      v_1166_0 <= 3'h0;
      v_1173_0 <= 3'h0;
      v_1180_0 <= 3'h0;
      v_1187_0 <= 3'h0;
      v_1194_0 <= 3'h0;
      v_1201_0 <= 3'h0;
      v_1208_0 <= 3'h0;
      v_1215_0 <= 3'h0;
      v_1222_0 <= 3'h0;
      v_1229_0 <= 3'h0;
      v_1236_0 <= 3'h0;
      v_1243_0 <= 3'h0;
      v_1250_0 <= 3'h0;
      v_1257_0 <= 3'h0;
      v_1264_0 <= 3'h0;
      v_1271_0 <= 3'h0;
      v_1278_0 <= 3'h0;
      v_1285_0 <= 3'h0;
      v_1292_0 <= 3'h0;
      v_1299_0 <= 3'h0;
      v_1306_0 <= 3'h0;
      v_1313_0 <= 3'h0;
      v_1320_0 <= 3'h0;
      v_1327_0 <= 3'h0;
      v_1334_0 <= 3'h0;
      v_1341_0 <= 3'h0;
      v_1348_0 <= 3'h0;
      v_1355_0 <= 3'h0;
      v_1362_0 <= 3'h0;
      v_1369_0 <= 3'h0;
      v_1376_0 <= 3'h0;
      v_1383_0 <= 3'h0;
      v_1390_0 <= 3'h0;
      v_1397_0 <= 3'h0;
      v_1404_0 <= 3'h0;
      v_1411_0 <= 3'h0;
      v_1418_0 <= 3'h0;
      v_1425_0 <= 3'h0;
      v_1432_0 <= 3'h0;
      v_1439_0 <= 3'h0;
      v_1446_0 <= 3'h0;
      v_1453_0 <= 3'h0;
      v_1460_0 <= 3'h0;
      v_1467_0 <= 3'h0;
      v_1474_0 <= 3'h0;
      v_1481_0 <= 3'h0;
      v_1488_0 <= 3'h0;
      v_1495_0 <= 3'h0;
      v_1502_0 <= 3'h0;
      v_1509_0 <= 3'h0;
      v_1516_0 <= 3'h0;
      v_1523_0 <= 3'h0;
      v_1530_0 <= 3'h0;
      v_1537_0 <= 3'h0;
      v_1544_0 <= 3'h0;
      v_1551_0 <= 3'h0;
      v_1558_0 <= 3'h0;
      v_1565_0 <= 3'h0;
      v_1572_0 <= 3'h0;
      v_1579_0 <= 3'h0;
      v_1586_0 <= 3'h0;
      v_1593_0 <= 3'h0;
      v_1600_0 <= 3'h0;
      v_1607_0 <= 3'h0;
      v_1614_0 <= 3'h0;
      v_1621_0 <= 3'h0;
      v_1628_0 <= 3'h0;
      v_1635_0 <= 3'h0;
      v_1642_0 <= 3'h0;
      v_1649_0 <= 3'h0;
      v_1656_0 <= 3'h0;
      v_1663_0 <= 3'h0;
      v_1670_0 <= 3'h0;
      v_1677_0 <= 3'h0;
      v_1684_0 <= 3'h0;
      v_1691_0 <= 3'h0;
      v_1698_0 <= 3'h0;
      v_1705_0 <= 3'h0;
      v_1712_0 <= 3'h0;
      v_1719_0 <= 3'h0;
      v_1726_0 <= 3'h0;
      v_1733_0 <= 3'h0;
      v_1740_0 <= 3'h0;
      v_1747_0 <= 3'h0;
      v_1754_0 <= 3'h0;
      v_1761_0 <= 3'h0;
      v_1768_0 <= 3'h0;
      v_1775_0 <= 3'h0;
      v_1782_0 <= 3'h0;
      v_1789_0 <= 3'h0;
      v_1796_0 <= 3'h0;
      v_1803_0 <= 3'h0;
      v_1810_0 <= 3'h0;
      v_1817_0 <= 3'h0;
      v_1824_0 <= 3'h0;
      v_1831_0 <= 3'h0;
      v_1838_0 <= 3'h0;
      v_1845_0 <= 3'h0;
      v_1852_0 <= 3'h0;
      v_1859_0 <= 3'h0;
      v_1866_0 <= 3'h0;
      v_1873_0 <= 3'h0;
      v_1880_0 <= 3'h0;
      v_1887_0 <= 3'h0;
      v_1894_0 <= 3'h0;
      v_1901_0 <= 3'h0;
      v_1908_0 <= 3'h0;
      v_1915_0 <= 3'h0;
      v_1922_0 <= 3'h0;
      v_1929_0 <= 3'h0;
      v_1936_0 <= 3'h0;
      v_1943_0 <= 3'h0;
      v_1950_0 <= 3'h0;
      v_1957_0 <= 3'h0;
      v_1964_0 <= 3'h0;
      v_1971_0 <= 3'h0;
      v_1978_0 <= 3'h0;
      v_1985_0 <= 3'h0;
      v_1992_0 <= 3'h0;
      v_1999_0 <= 3'h0;
      v_2006_0 <= 3'h0;
      v_2013_0 <= 3'h0;
      v_2020_0 <= 3'h0;
      v_2027_0 <= 3'h0;
      v_2034_0 <= 3'h0;
      v_2041_0 <= 3'h0;
      v_2048_0 <= 3'h0;
      v_2055_0 <= 3'h0;
      v_2062_0 <= 3'h0;
      v_2069_0 <= 3'h0;
      v_2076_0 <= 3'h0;
      v_2083_0 <= 3'h0;
      v_2090_0 <= 3'h0;
      v_2097_0 <= 3'h0;
      v_2104_0 <= 3'h0;
      v_2111_0 <= 3'h0;
      v_2118_0 <= 3'h0;
      v_2125_0 <= 3'h0;
      v_2132_0 <= 3'h0;
      v_2139_0 <= 3'h0;
      v_2146_0 <= 3'h0;
      v_2153_0 <= 3'h0;
      v_2160_0 <= 3'h0;
      v_2167_0 <= 3'h0;
      v_2174_0 <= 3'h0;
      v_2181_0 <= 3'h0;
      v_2188_0 <= 3'h0;
      v_2195_0 <= 3'h0;
      v_2202_0 <= 3'h0;
      v_2209_0 <= 3'h0;
      v_2216_0 <= 3'h0;
      v_2223_0 <= 3'h0;
      v_2230_0 <= 3'h0;
      v_2237_0 <= 3'h0;
      v_2244_0 <= 3'h0;
      v_2251_0 <= 3'h0;
      v_2258_0 <= 3'h0;
      v_2265_0 <= 3'h0;
      v_2272_0 <= 3'h0;
      v_2279_0 <= 3'h0;
      v_2286_0 <= 3'h0;
      v_2293_0 <= 3'h0;
      v_2300_0 <= 3'h0;
      v_2307_0 <= 3'h0;
      v_2314_0 <= 3'h0;
      v_2321_0 <= 3'h0;
      v_2328_0 <= 3'h0;
      v_2335_0 <= 3'h0;
      v_2342_0 <= 3'h0;
      v_2349_0 <= 3'h0;
      v_2356_0 <= 3'h0;
      v_2363_0 <= 3'h0;
      v_2370_0 <= 3'h0;
      v_2377_0 <= 3'h0;
      v_2384_0 <= 3'h0;
      v_2391_0 <= 3'h0;
      v_2398_0 <= 3'h0;
      v_2405_0 <= 3'h0;
      v_2412_0 <= 3'h0;
      v_2419_0 <= 3'h0;
      v_2426_0 <= 3'h0;
      v_2433_0 <= 3'h0;
      v_2440_0 <= 3'h0;
      v_2447_0 <= 3'h0;
      v_2454_0 <= 3'h0;
      v_2461_0 <= 3'h0;
      v_2468_0 <= 3'h0;
      v_2475_0 <= 3'h0;
      v_2482_0 <= 3'h0;
      v_2489_0 <= 3'h0;
      v_2496_0 <= 3'h0;
      v_2503_0 <= 3'h0;
      v_2510_0 <= 3'h0;
      v_2517_0 <= 3'h0;
      v_2524_0 <= 3'h0;
      v_2531_0 <= 3'h0;
      v_2538_0 <= 3'h0;
      v_2545_0 <= 3'h0;
      v_2552_0 <= 3'h0;
      v_2559_0 <= 3'h0;
      v_2566_0 <= 3'h0;
      v_2573_0 <= 3'h0;
      v_2580_0 <= 3'h0;
      v_2587_0 <= 3'h0;
      v_2594_0 <= 3'h0;
      v_2601_0 <= 3'h0;
      v_2608_0 <= 3'h0;
      v_2615_0 <= 3'h0;
      v_2622_0 <= 3'h0;
      v_2629_0 <= 3'h0;
      v_2636_0 <= 3'h0;
      v_2643_0 <= 3'h0;
      v_2650_0 <= 3'h0;
      v_2657_0 <= 3'h0;
      v_2664_0 <= 3'h0;
      v_2671_0 <= 3'h0;
      v_2678_0 <= 3'h0;
      v_2685_0 <= 3'h0;
      v_2692_0 <= 3'h0;
      v_2699_0 <= 3'h0;
      v_2706_0 <= 3'h0;
      v_2713_0 <= 3'h0;
      v_2720_0 <= 3'h0;
      v_2727_0 <= 3'h0;
      v_2734_0 <= 3'h0;
      v_2741_0 <= 3'h0;
      v_2748_0 <= 3'h0;
      v_2755_0 <= 3'h0;
      v_2762_0 <= 3'h0;
      v_2769_0 <= 3'h0;
      v_2776_0 <= 3'h0;
      v_2783_0 <= 3'h0;
      v_2790_0 <= 3'h0;
      v_2797_0 <= 3'h0;
      v_2804_0 <= 3'h0;
      v_2811_0 <= 3'h0;
      v_2818_0 <= 3'h0;
      v_2825_0 <= 3'h0;
      v_2832_0 <= 3'h0;
      v_2839_0 <= 3'h0;
      v_2846_0 <= 3'h0;
      v_2853_0 <= 3'h0;
      v_2860_0 <= 3'h0;
      v_2867_0 <= 3'h0;
      v_2874_0 <= 3'h0;
      v_2881_0 <= 3'h0;
      v_2888_0 <= 3'h0;
      v_2895_0 <= 3'h0;
      v_2902_0 <= 3'h0;
      v_2909_0 <= 3'h0;
      v_2916_0 <= 3'h0;
      v_2923_0 <= 3'h0;
      v_2930_0 <= 3'h0;
      v_2937_0 <= 3'h0;
      v_2944_0 <= 3'h0;
      v_2951_0 <= 3'h0;
      v_2958_0 <= 3'h0;
      v_2965_0 <= 3'h0;
      v_2972_0 <= 3'h0;
      v_2979_0 <= 3'h0;
      v_2986_0 <= 3'h0;
      v_2993_0 <= 3'h0;
      v_3000_0 <= 3'h0;
      v_3007_0 <= 3'h0;
      v_3014_0 <= 3'h0;
      v_3021_0 <= 3'h0;
      v_3028_0 <= 3'h0;
      v_3035_0 <= 3'h0;
      v_3042_0 <= 3'h0;
      v_3049_0 <= 3'h0;
      v_3056_0 <= 3'h0;
      v_3063_0 <= 3'h0;
      v_3070_0 <= 3'h0;
      v_3077_0 <= 3'h0;
      v_3084_0 <= 3'h0;
      v_3091_0 <= 3'h0;
      v_3098_0 <= 3'h0;
      v_3105_0 <= 3'h0;
      v_3112_0 <= 3'h0;
      v_3119_0 <= 3'h0;
      v_3126_0 <= 3'h0;
      v_3133_0 <= 3'h0;
      v_3140_0 <= 3'h0;
      v_3147_0 <= 3'h0;
      v_3154_0 <= 3'h0;
      v_3161_0 <= 3'h0;
      v_3168_0 <= 3'h0;
      v_3175_0 <= 3'h0;
      v_3182_0 <= 3'h0;
      v_3189_0 <= 3'h0;
      v_3196_0 <= 3'h0;
      v_3203_0 <= 3'h0;
      v_3210_0 <= 3'h0;
      v_3217_0 <= 3'h0;
      v_3224_0 <= 3'h0;
      v_3231_0 <= 3'h0;
      v_3238_0 <= 3'h0;
      v_3245_0 <= 3'h0;
      v_3252_0 <= 3'h0;
      v_3259_0 <= 3'h0;
      v_3266_0 <= 3'h0;
      v_3273_0 <= 3'h0;
      v_3280_0 <= 3'h0;
      v_3287_0 <= 3'h0;
      v_3294_0 <= 3'h0;
      v_3301_0 <= 3'h0;
      v_3308_0 <= 3'h0;
      v_3315_0 <= 3'h0;
      v_3322_0 <= 3'h0;
      v_3329_0 <= 3'h0;
      v_3336_0 <= 3'h0;
      v_3343_0 <= 3'h0;
      v_3350_0 <= 3'h0;
      v_3357_0 <= 3'h0;
      v_3364_0 <= 3'h0;
      v_3371_0 <= 3'h0;
      v_3378_0 <= 3'h0;
      v_3385_0 <= 3'h0;
      v_3392_0 <= 3'h0;
      v_3399_0 <= 3'h0;
      v_3406_0 <= 3'h0;
      v_3413_0 <= 3'h0;
      v_3420_0 <= 3'h0;
      v_3427_0 <= 3'h0;
      v_3434_0 <= 3'h0;
      v_3441_0 <= 3'h0;
      v_3448_0 <= 3'h0;
      v_3455_0 <= 3'h0;
      v_3462_0 <= 3'h0;
      v_3469_0 <= 3'h0;
      v_3476_0 <= 3'h0;
      v_3483_0 <= 3'h0;
      v_3490_0 <= 3'h0;
      v_3497_0 <= 3'h0;
      v_3504_0 <= 3'h0;
      v_3511_0 <= 3'h0;
      v_3518_0 <= 3'h0;
      v_3525_0 <= 3'h0;
      v_3532_0 <= 3'h0;
      v_3539_0 <= 3'h0;
      v_3546_0 <= 3'h0;
      v_3553_0 <= 3'h0;
      v_3560_0 <= 3'h0;
      v_3567_0 <= 3'h0;
      v_3574_0 <= 3'h0;
      v_3581_0 <= 3'h0;
      v_3588_0 <= 3'h0;
      v_3595_0 <= 3'h0;
      v_3602_0 <= 3'h0;
      v_3609_0 <= 3'h0;
      v_3616_0 <= 3'h0;
      v_3623_0 <= 3'h0;
      v_3630_0 <= 3'h0;
      v_3637_0 <= 3'h0;
      v_3644_0 <= 3'h0;
      v_3651_0 <= 3'h0;
      v_3658_0 <= 3'h0;
      v_3665_0 <= 3'h0;
      v_3672_0 <= 3'h0;
      v_3679_0 <= 3'h0;
      v_3686_0 <= 3'h0;
      v_3693_0 <= 3'h0;
      v_3700_0 <= 3'h0;
      v_3707_0 <= 3'h0;
      v_3714_0 <= 3'h0;
      v_3721_0 <= 3'h0;
      v_3728_0 <= 3'h0;
      v_3735_0 <= 3'h0;
      v_3742_0 <= 3'h0;
      v_3749_0 <= 3'h0;
      v_3756_0 <= 3'h0;
      v_3763_0 <= 3'h0;
      v_3770_0 <= 3'h0;
      v_3777_0 <= 3'h0;
      v_3784_0 <= 3'h0;
      v_3791_0 <= 3'h0;
      v_3798_0 <= 3'h0;
      v_3805_0 <= 3'h0;
      v_3812_0 <= 3'h0;
      v_3819_0 <= 3'h0;
      v_3826_0 <= 3'h0;
      v_3833_0 <= 3'h0;
      v_3840_0 <= 3'h0;
      v_3847_0 <= 3'h0;
      v_3854_0 <= 3'h0;
      v_3861_0 <= 3'h0;
      v_3868_0 <= 3'h0;
      v_3875_0 <= 3'h0;
      v_3882_0 <= 3'h0;
      v_3889_0 <= 3'h0;
      v_3896_0 <= 3'h0;
      v_3903_0 <= 3'h0;
      v_3910_0 <= 3'h0;
      v_3917_0 <= 3'h0;
      v_3924_0 <= 3'h0;
      v_3931_0 <= 3'h0;
      v_3938_0 <= 3'h0;
      v_3945_0 <= 3'h0;
      v_3952_0 <= 3'h0;
      v_3959_0 <= 3'h0;
      v_3966_0 <= 3'h0;
      v_3973_0 <= 3'h0;
      v_3980_0 <= 3'h0;
      v_3987_0 <= 3'h0;
      v_3994_0 <= 3'h0;
      v_4001_0 <= 3'h0;
      v_4008_0 <= 3'h0;
      v_4015_0 <= 3'h0;
      v_4022_0 <= 3'h0;
      v_4029_0 <= 3'h0;
      v_4036_0 <= 3'h0;
      v_4043_0 <= 3'h0;
      v_4050_0 <= 3'h0;
      v_4057_0 <= 3'h0;
      v_4064_0 <= 3'h0;
      v_4071_0 <= 3'h0;
      v_4078_0 <= 3'h0;
      v_4085_0 <= 3'h0;
      v_4092_0 <= 3'h0;
      v_4099_0 <= 3'h0;
      v_4106_0 <= 3'h0;
      v_4113_0 <= 3'h0;
      v_4120_0 <= 3'h0;
      v_4127_0 <= 3'h0;
      v_4134_0 <= 3'h0;
      v_4141_0 <= 3'h0;
      v_4148_0 <= 3'h0;
      v_4155_0 <= 3'h0;
      v_4162_0 <= 3'h0;
      v_4169_0 <= 3'h0;
      v_4176_0 <= 3'h0;
      v_4183_0 <= 3'h0;
      v_4190_0 <= 3'h0;
      v_4197_0 <= 3'h0;
      v_4204_0 <= 3'h0;
      v_4211_0 <= 3'h0;
      v_4218_0 <= 3'h0;
      v_4225_0 <= 3'h0;
      v_4232_0 <= 3'h0;
      v_4239_0 <= 3'h0;
      v_4246_0 <= 3'h0;
      v_4253_0 <= 3'h0;
      v_4260_0 <= 3'h0;
      v_4267_0 <= 3'h0;
      v_4274_0 <= 3'h0;
      v_4281_0 <= 3'h0;
      v_4288_0 <= 3'h0;
      v_4295_0 <= 3'h0;
      v_4302_0 <= 3'h0;
      v_4309_0 <= 3'h0;
      v_4316_0 <= 3'h0;
      v_4323_0 <= 3'h0;
      v_4330_0 <= 3'h0;
      v_4337_0 <= 3'h0;
      v_4344_0 <= 3'h0;
      v_4351_0 <= 3'h0;
      v_4358_0 <= 3'h0;
      v_4365_0 <= 3'h0;
      v_4372_0 <= 3'h0;
      v_4379_0 <= 3'h0;
      v_4386_0 <= 3'h0;
      v_4393_0 <= 3'h0;
      v_4400_0 <= 3'h0;
      v_4407_0 <= 3'h0;
      v_4414_0 <= 3'h0;
      v_4421_0 <= 3'h0;
      v_4428_0 <= 3'h0;
      v_4435_0 <= 3'h0;
      v_4442_0 <= 3'h0;
      v_4449_0 <= 3'h0;
      v_4456_0 <= 3'h0;
      v_4463_0 <= 3'h0;
      v_4470_0 <= 3'h0;
      v_4477_0 <= 3'h0;
      v_4484_0 <= 3'h0;
      v_4491_0 <= 3'h0;
      v_4498_0 <= 3'h0;
      v_4505_0 <= 3'h0;
      v_4512_0 <= 3'h0;
      v_4519_0 <= 3'h0;
      v_4526_0 <= 3'h0;
      v_4533_0 <= 3'h0;
      v_4540_0 <= 3'h0;
      v_4547_0 <= 3'h0;
      v_4554_0 <= 3'h0;
      v_4561_0 <= 3'h0;
      v_4568_0 <= 3'h0;
      v_4575_0 <= 3'h0;
      v_4582_0 <= 3'h0;
      v_4589_0 <= 3'h0;
      v_4596_0 <= 3'h0;
      v_4603_0 <= 3'h0;
      v_4610_0 <= 3'h0;
      v_4617_0 <= 3'h0;
      v_4624_0 <= 3'h0;
      v_4631_0 <= 3'h0;
      v_4638_0 <= 3'h0;
      v_4645_0 <= 3'h0;
      v_4652_0 <= 3'h0;
      v_4659_0 <= 3'h0;
      v_4666_0 <= 3'h0;
      v_4673_0 <= 3'h0;
      v_4680_0 <= 3'h0;
      v_4687_0 <= 3'h0;
      v_4694_0 <= 3'h0;
      v_4701_0 <= 3'h0;
      v_4708_0 <= 3'h0;
      v_4715_0 <= 3'h0;
      v_4722_0 <= 3'h0;
      v_4729_0 <= 3'h0;
      v_4736_0 <= 3'h0;
      v_4743_0 <= 3'h0;
      v_4750_0 <= 3'h0;
      v_4757_0 <= 3'h0;
      v_4764_0 <= 3'h0;
      v_4771_0 <= 3'h0;
      v_4778_0 <= 3'h0;
      v_4785_0 <= 3'h0;
      v_4792_0 <= 3'h0;
      v_4799_0 <= 3'h0;
      v_4806_0 <= 3'h0;
      v_4813_0 <= 3'h0;
      v_4820_0 <= 3'h0;
      v_4827_0 <= 3'h0;
      v_4834_0 <= 3'h0;
      v_4841_0 <= 3'h0;
      v_4848_0 <= 3'h0;
      v_4855_0 <= 3'h0;
      v_4862_0 <= 3'h0;
      v_4869_0 <= 3'h0;
      v_4876_0 <= 3'h0;
      v_4883_0 <= 3'h0;
      v_4890_0 <= 3'h0;
      v_4897_0 <= 3'h0;
      v_4904_0 <= 3'h0;
      v_4911_0 <= 3'h0;
      v_4918_0 <= 3'h0;
      v_4925_0 <= 3'h0;
      v_4932_0 <= 3'h0;
      v_4939_0 <= 3'h0;
      v_4946_0 <= 3'h0;
      v_4953_0 <= 3'h0;
      v_4960_0 <= 3'h0;
      v_4967_0 <= 3'h0;
      v_4974_0 <= 3'h0;
      v_4981_0 <= 3'h0;
      v_4988_0 <= 3'h0;
      v_4995_0 <= 3'h0;
      v_5002_0 <= 3'h0;
      v_5009_0 <= 3'h0;
      v_5016_0 <= 3'h0;
      v_5023_0 <= 3'h0;
      v_5030_0 <= 3'h0;
      v_5037_0 <= 3'h0;
      v_5044_0 <= 3'h0;
      v_5051_0 <= 3'h0;
      v_5058_0 <= 3'h0;
      v_5065_0 <= 3'h0;
      v_5072_0 <= 3'h0;
      v_5079_0 <= 3'h0;
      v_5086_0 <= 3'h0;
      v_5093_0 <= 3'h0;
      v_5100_0 <= 3'h0;
      v_5107_0 <= 3'h0;
      v_5114_0 <= 3'h0;
      v_5121_0 <= 3'h0;
      v_5128_0 <= 3'h0;
      v_5135_0 <= 3'h0;
      v_5142_0 <= 3'h0;
      v_5149_0 <= 3'h0;
      v_5156_0 <= 3'h0;
      v_5163_0 <= 3'h0;
      v_5170_0 <= 3'h0;
      v_5177_0 <= 3'h0;
      v_5184_0 <= 3'h0;
      v_5191_0 <= 3'h0;
      v_5198_0 <= 3'h0;
      v_5205_0 <= 3'h0;
      v_5212_0 <= 3'h0;
      v_5219_0 <= 3'h0;
      v_5226_0 <= 3'h0;
      v_5233_0 <= 3'h0;
      v_5240_0 <= 3'h0;
      v_5247_0 <= 3'h0;
      v_5254_0 <= 3'h0;
      v_5261_0 <= 3'h0;
      v_5268_0 <= 3'h0;
      v_5275_0 <= 3'h0;
      v_5282_0 <= 3'h0;
      v_5289_0 <= 3'h0;
      v_5296_0 <= 3'h0;
      v_5303_0 <= 3'h0;
      v_5310_0 <= 3'h0;
      v_5317_0 <= 3'h0;
      v_5324_0 <= 3'h0;
      v_5331_0 <= 3'h0;
      v_5338_0 <= 3'h0;
      v_5345_0 <= 3'h0;
      v_5352_0 <= 3'h0;
      v_5359_0 <= 3'h0;
      v_5366_0 <= 3'h0;
      v_5373_0 <= 3'h0;
      v_5380_0 <= 3'h0;
      v_5387_0 <= 3'h0;
      v_5394_0 <= 3'h0;
      v_5401_0 <= 3'h0;
      v_5408_0 <= 3'h0;
      v_5415_0 <= 3'h0;
      v_5422_0 <= 3'h0;
      v_5429_0 <= 3'h0;
      v_5436_0 <= 3'h0;
      v_5443_0 <= 3'h0;
      v_5450_0 <= 3'h0;
      v_5457_0 <= 3'h0;
      v_5464_0 <= 3'h0;
      v_5471_0 <= 3'h0;
      v_5478_0 <= 3'h0;
      v_5485_0 <= 3'h0;
      v_5492_0 <= 3'h0;
      v_5499_0 <= 3'h0;
      v_5506_0 <= 3'h0;
      v_5513_0 <= 3'h0;
      v_5520_0 <= 3'h0;
      v_5527_0 <= 3'h0;
      v_5534_0 <= 3'h0;
      v_5541_0 <= 3'h0;
      v_5548_0 <= 3'h0;
      v_5555_0 <= 3'h0;
      v_5562_0 <= 3'h0;
      v_5569_0 <= 3'h0;
      v_5576_0 <= 3'h0;
      v_5583_0 <= 3'h0;
      v_5590_0 <= 3'h0;
      v_5597_0 <= 3'h0;
      v_5604_0 <= 3'h0;
      v_5611_0 <= 3'h0;
      v_5618_0 <= 3'h0;
      v_5625_0 <= 3'h0;
      v_5632_0 <= 3'h0;
      v_5639_0 <= 3'h0;
      v_5646_0 <= 3'h0;
      v_5653_0 <= 3'h0;
      v_5660_0 <= 3'h0;
      v_5667_0 <= 3'h0;
      v_5674_0 <= 3'h0;
      v_5681_0 <= 3'h0;
      v_5688_0 <= 3'h0;
      v_5695_0 <= 3'h0;
      v_5702_0 <= 3'h0;
      v_5709_0 <= 3'h0;
      v_5716_0 <= 3'h0;
      v_5723_0 <= 3'h0;
      v_5730_0 <= 3'h0;
      v_5737_0 <= 3'h0;
      v_5744_0 <= 3'h0;
      v_5751_0 <= 3'h0;
      v_5758_0 <= 3'h0;
      v_5765_0 <= 3'h0;
      v_5772_0 <= 3'h0;
      v_5779_0 <= 3'h0;
      v_5786_0 <= 3'h0;
      v_5793_0 <= 3'h0;
      v_5800_0 <= 3'h0;
      v_5807_0 <= 3'h0;
      v_5814_0 <= 3'h0;
      v_5821_0 <= 3'h0;
      v_5828_0 <= 3'h0;
      v_5835_0 <= 3'h0;
      v_5842_0 <= 3'h0;
      v_5849_0 <= 3'h0;
      v_5856_0 <= 3'h0;
      v_5863_0 <= 3'h0;
      v_5870_0 <= 3'h0;
      v_5877_0 <= 3'h0;
      v_5884_0 <= 3'h0;
      v_5891_0 <= 3'h0;
      v_5898_0 <= 3'h0;
      v_5905_0 <= 3'h0;
      v_5912_0 <= 3'h0;
      v_5919_0 <= 3'h0;
      v_5926_0 <= 3'h0;
      v_5933_0 <= 3'h0;
      v_5940_0 <= 3'h0;
      v_5947_0 <= 3'h0;
      v_5954_0 <= 3'h0;
      v_5961_0 <= 3'h0;
      v_5968_0 <= 3'h0;
      v_5975_0 <= 3'h0;
      v_5982_0 <= 3'h0;
      v_5989_0 <= 3'h0;
      v_5996_0 <= 3'h0;
      v_6003_0 <= 3'h0;
      v_6010_0 <= 3'h0;
      v_6017_0 <= 3'h0;
      v_6024_0 <= 3'h0;
      v_6031_0 <= 3'h0;
      v_6038_0 <= 3'h0;
      v_6045_0 <= 3'h0;
      v_6052_0 <= 3'h0;
      v_6059_0 <= 3'h0;
      v_6066_0 <= 3'h0;
      v_6073_0 <= 3'h0;
      v_6080_0 <= 3'h0;
      v_6087_0 <= 3'h0;
      v_6094_0 <= 3'h0;
      v_6101_0 <= 3'h0;
      v_6108_0 <= 3'h0;
      v_6115_0 <= 3'h0;
      v_6122_0 <= 3'h0;
      v_6129_0 <= 3'h0;
      v_6136_0 <= 3'h0;
      v_6143_0 <= 3'h0;
      v_6150_0 <= 3'h0;
      v_6157_0 <= 3'h0;
      v_6164_0 <= 3'h0;
      v_6171_0 <= 3'h0;
      v_6178_0 <= 3'h0;
      v_6185_0 <= 3'h0;
      v_6192_0 <= 3'h0;
      v_6199_0 <= 3'h0;
      v_6206_0 <= 3'h0;
      v_6213_0 <= 3'h0;
      v_6220_0 <= 3'h0;
      v_6227_0 <= 3'h0;
      v_6234_0 <= 3'h0;
      v_6241_0 <= 3'h0;
      v_6248_0 <= 3'h0;
      v_6255_0 <= 3'h0;
      v_6262_0 <= 3'h0;
      v_6269_0 <= 3'h0;
      v_6276_0 <= 3'h0;
      v_6283_0 <= 3'h0;
      v_6290_0 <= 3'h0;
      v_6297_0 <= 3'h0;
      v_6304_0 <= 3'h0;
      v_6311_0 <= 3'h0;
      v_6318_0 <= 3'h0;
      v_6325_0 <= 3'h0;
      v_6332_0 <= 3'h0;
      v_6339_0 <= 3'h0;
      v_6346_0 <= 3'h0;
      v_6353_0 <= 3'h0;
      v_6360_0 <= 3'h0;
      v_6367_0 <= 3'h0;
      v_6374_0 <= 3'h0;
      v_6381_0 <= 3'h0;
      v_6388_0 <= 3'h0;
      v_6395_0 <= 3'h0;
      v_6402_0 <= 3'h0;
      v_6409_0 <= 3'h0;
      v_6416_0 <= 3'h0;
      v_6423_0 <= 3'h0;
      v_6430_0 <= 3'h0;
      v_6437_0 <= 3'h0;
      v_6444_0 <= 3'h0;
      v_6451_0 <= 3'h0;
      v_6458_0 <= 3'h0;
      v_6465_0 <= 3'h0;
      v_6472_0 <= 3'h0;
      v_6479_0 <= 3'h0;
      v_6486_0 <= 3'h0;
      v_6493_0 <= 3'h0;
      v_6500_0 <= 3'h0;
      v_6507_0 <= 3'h0;
      v_6514_0 <= 3'h0;
      v_6521_0 <= 3'h0;
      v_6528_0 <= 3'h0;
      v_6535_0 <= 3'h0;
      v_6542_0 <= 3'h0;
      v_6549_0 <= 3'h0;
      v_6556_0 <= 3'h0;
      v_6563_0 <= 3'h0;
      v_6570_0 <= 3'h0;
      v_6577_0 <= 3'h0;
      v_6584_0 <= 3'h0;
      v_6591_0 <= 3'h0;
      v_6598_0 <= 3'h0;
      v_6605_0 <= 3'h0;
      v_6612_0 <= 3'h0;
      v_6619_0 <= 3'h0;
      v_6626_0 <= 3'h0;
      v_6633_0 <= 3'h0;
      v_6640_0 <= 3'h0;
      v_6647_0 <= 3'h0;
      v_6654_0 <= 3'h0;
      v_6661_0 <= 3'h0;
      v_6668_0 <= 3'h0;
      v_6675_0 <= 3'h0;
      v_6682_0 <= 3'h0;
      v_6689_0 <= 3'h0;
      v_6696_0 <= 3'h0;
      v_6703_0 <= 3'h0;
      v_6710_0 <= 3'h0;
      v_6717_0 <= 3'h0;
      v_6724_0 <= 3'h0;
      v_6731_0 <= 3'h0;
      v_6738_0 <= 3'h0;
      v_6745_0 <= 3'h0;
      v_6752_0 <= 3'h0;
      v_6759_0 <= 3'h0;
      v_6766_0 <= 3'h0;
      v_6773_0 <= 3'h0;
      v_6780_0 <= 3'h0;
      v_6787_0 <= 3'h0;
      v_6794_0 <= 3'h0;
      v_6801_0 <= 3'h0;
      v_6808_0 <= 3'h0;
      v_6815_0 <= 3'h0;
      v_6822_0 <= 3'h0;
      v_6829_0 <= 3'h0;
      v_6836_0 <= 3'h0;
      v_6843_0 <= 3'h0;
      v_6850_0 <= 3'h0;
      v_6857_0 <= 3'h0;
      v_6864_0 <= 3'h0;
      v_6871_0 <= 3'h0;
      v_6878_0 <= 3'h0;
      v_6885_0 <= 3'h0;
      v_6892_0 <= 3'h0;
      v_6899_0 <= 3'h0;
      v_6906_0 <= 3'h0;
      v_6913_0 <= 3'h0;
      v_6920_0 <= 3'h0;
      v_6927_0 <= 3'h0;
      v_6934_0 <= 3'h0;
      v_6941_0 <= 3'h0;
      v_6948_0 <= 3'h0;
      v_6955_0 <= 3'h0;
      v_6962_0 <= 3'h0;
      v_6969_0 <= 3'h0;
      v_6976_0 <= 3'h0;
      v_6983_0 <= 3'h0;
      v_6990_0 <= 3'h0;
      v_6997_0 <= 3'h0;
      v_7004_0 <= 3'h0;
      v_7011_0 <= 3'h0;
      v_7018_0 <= 3'h0;
      v_7025_0 <= 3'h0;
      v_7032_0 <= 3'h0;
      v_7039_0 <= 3'h0;
      v_7046_0 <= 3'h0;
      v_7053_0 <= 3'h0;
      v_7060_0 <= 3'h0;
      v_7067_0 <= 3'h0;
      v_7074_0 <= 3'h0;
      v_7081_0 <= 3'h0;
      v_7088_0 <= 3'h0;
      v_7095_0 <= 3'h0;
      v_7102_0 <= 3'h0;
      v_7109_0 <= 3'h0;
      v_7116_0 <= 3'h0;
      v_7123_0 <= 3'h0;
      v_7130_0 <= 3'h0;
      v_7137_0 <= 3'h0;
      v_7144_0 <= 3'h0;
      v_7151_0 <= 3'h0;
      v_7158_0 <= 3'h0;
      v_7165_0 <= 3'h0;
      v_7172_0 <= 3'h0;
      v_7179_0 <= 3'h0;
      v_7186_0 <= 3'h0;
      v_7193_0 <= 3'h0;
      v_7200_0 <= 3'h0;
      v_7207_0 <= 3'h0;
      v_7214_0 <= 3'h0;
      v_7221_0 <= 3'h0;
      v_7228_0 <= 3'h0;
      v_7235_0 <= 3'h0;
      v_7242_0 <= 3'h0;
      v_7249_0 <= 3'h0;
      v_7256_0 <= 3'h0;
      v_7263_0 <= 3'h0;
      v_7270_0 <= 3'h0;
      v_7277_0 <= 3'h0;
      v_7284_0 <= 3'h0;
      v_7291_0 <= 3'h0;
      v_7298_0 <= 3'h0;
      v_7305_0 <= 3'h0;
      v_7312_0 <= 3'h0;
      v_7319_0 <= 3'h0;
      v_7326_0 <= 3'h0;
      v_7333_0 <= 3'h0;
      v_7340_0 <= 3'h0;
      v_7347_0 <= 3'h0;
      v_7354_0 <= 3'h0;
      v_7361_0 <= 3'h0;
      v_7368_0 <= 3'h0;
      v_7375_0 <= 3'h0;
      v_7382_0 <= 3'h0;
      v_7389_0 <= 3'h0;
      v_7396_0 <= 3'h0;
      v_7403_0 <= 3'h0;
      v_7410_0 <= 3'h0;
      v_7417_0 <= 3'h0;
      v_7424_0 <= 3'h0;
      v_7431_0 <= 3'h0;
      v_7438_0 <= 3'h0;
      v_7445_0 <= 3'h0;
      v_7452_0 <= 3'h0;
      v_7459_0 <= 3'h0;
      v_7466_0 <= 3'h0;
      v_7473_0 <= 3'h0;
      v_7480_0 <= 3'h0;
      v_7487_0 <= 3'h0;
      v_7494_0 <= 3'h0;
      v_7501_0 <= 3'h0;
      v_7508_0 <= 3'h0;
      v_7515_0 <= 3'h0;
      v_7522_0 <= 3'h0;
      v_7529_0 <= 3'h0;
      v_7536_0 <= 3'h0;
      v_7543_0 <= 3'h0;
      v_7550_0 <= 3'h0;
      v_7557_0 <= 3'h0;
      v_7564_0 <= 3'h0;
      v_7571_0 <= 3'h0;
      v_7578_0 <= 3'h0;
      v_7585_0 <= 3'h0;
      v_7592_0 <= 3'h0;
      v_7599_0 <= 3'h0;
      v_7606_0 <= 3'h0;
      v_7613_0 <= 3'h0;
      v_7620_0 <= 3'h0;
      v_7627_0 <= 3'h0;
      v_7634_0 <= 3'h0;
      v_7641_0 <= 3'h0;
      v_7648_0 <= 3'h0;
      v_7655_0 <= 3'h0;
      v_7662_0 <= 3'h0;
      v_7669_0 <= 3'h0;
      v_7676_0 <= 3'h0;
      v_7683_0 <= 3'h0;
      v_7690_0 <= 3'h0;
      v_7697_0 <= 3'h0;
      v_7704_0 <= 3'h0;
      v_7711_0 <= 3'h0;
      v_7718_0 <= 3'h0;
      v_7725_0 <= 3'h0;
      v_7732_0 <= 3'h0;
      v_7739_0 <= 3'h0;
      v_7746_0 <= 3'h0;
      v_7753_0 <= 3'h0;
      v_7760_0 <= 3'h0;
      v_7767_0 <= 3'h0;
      v_7774_0 <= 3'h0;
      v_7781_0 <= 3'h0;
      v_7788_0 <= 3'h0;
      v_7795_0 <= 3'h0;
      v_7802_0 <= 3'h0;
      v_7809_0 <= 3'h0;
      v_7816_0 <= 3'h0;
      v_7823_0 <= 3'h0;
      v_7830_0 <= 3'h0;
      v_7837_0 <= 3'h0;
      v_7844_0 <= 3'h0;
      v_7851_0 <= 3'h0;
      v_11948_0 <= 3'h0;
      v_11960_0 <= 1'h0;
      v_11961_0 <= 1'h0;
      v_11965_0 <= 10'h0;
      v_11989_0 <= 10'h0;
      v_11993_0 <= 10'h0;
      v_12002_0 <= 3'h0;
      v_12065_0 <= 1'h1;
      v_12078_0 <= 1'h0;
      v_12086_0 <= 16'h0;
      v_12090_0 <= 1'h0;
      v_12092_0 <= 1'h0;
      v_12099_0 <= 1'h1;
      v_12109_0 <= 5'h0;
      v_12110_0 <= 5'h0;
      v_12156_0 <= 16'h0;
      v_12170_0 <= 1'h0;
      v_12171_0 <= 1'h0;
      v_12173_0 <= 5'h0;
      v_12178_0 <= 5'h0;
      v_12183_0 <= 16'h0;
      v_12226_0 <= 16'h0;
      v_12288_0 <= 1'h0;
      v_12294_0 <= 32'h0;
      v_12334_0 <= 1'h0;
      v_12345_0 <= 1'h0;
      v_12356_0 <= 8'h0;
      v_12358_0 <= 8'h0;
    end else begin
      if (v_1_0 == 1) $write ("Push", " ");
      if (v_4_0 == 1) v_3_0 <= 1'h1;
      if (v_13_0 == 1) v_12_0 <= v_12085_0;
      if (v_19_0 == 1) v_18_0 <= 1'h1;
      if (v_24_0 == 1) v_23_0 <= v_676_0;
      if (v_35_0 == 1) v_34_0 <= v_579_0;
      if (v_41_0 == 1) v_40_0 <= v_568_0;
      if (v_13_0 == 1) v_52_0 <= v_53_0;
      if (v_55_0 == 1) v_54_0 <= v_190_0;
      if (v_55_0 == 1) v_58_0 <= v_59_0;
      if (v_61_0 == 1) v_60_0 <= v_174_0;
      if (v_68_0 == 1) v_67_0 <= v_168_0;
      if (1'h1 == 1) v_77_0 <= v_71_0;
      if (_act_79_0 == 1) v_78_0 <= v_162_0;
      if (v_92_0 == 1) v_91_0 <= v_114_0;
      if (v_98_0 == 1) v_97_0 <= v_105_0;
      if (v_192_0 == 1) v_191_0 <= v_200_0;
      v_205_0 <= 1'h1;
      v_206_0 <= _act_79_0;
      v_208_0 <= v_209_0;
      v_213_0 <= v_214_0;
      v_218_0 <= v_219_0;
      if (v_272_0 == 1) v_271_0 <= v_301_0;
      if (v_13_0 == 1) v_330_0 <= v_331_0;
      if (v_333_0 == 1) v_332_0 <= v_433_0;
      if (v_333_0 == 1) v_336_0 <= v_337_0;
      if (v_339_0 == 1) v_338_0 <= v_417_0;
      if (v_346_0 == 1) v_345_0 <= v_411_0;
      if (1'h1 == 1) v_355_0 <= v_349_0;
      if (_act_357_0 == 1) v_356_0 <= v_405_0;
      if (v_435_0 == 1) v_434_0 <= v_443_0;
      v_448_0 <= 1'h1;
      v_449_0 <= _act_357_0;
      v_451_0 <= v_452_0;
      v_456_0 <= v_457_0;
      v_461_0 <= v_462_0;
      if (v_515_0 == 1) v_514_0 <= v_544_0;
      if (v_13_0 == 1) v_578_0 <= v_12_0;
      if (v_598_0 == 1) v_597_0 <= v_657_0;
      v_615_0 <= v_616_0;
      if (v_617_0 == 1) v_616_0 <= v_649_0;
      if (v_621_0 == 1) v_620_0 <= v_638_0;
      v_642_0 <= v_615_0;
      if (v_691_0 == 1) v_690_0 <= v_694_0;
      if (v_698_0 == 1) v_697_0 <= v_701_0;
      if (v_705_0 == 1) v_704_0 <= v_708_0;
      if (v_712_0 == 1) v_711_0 <= v_715_0;
      if (v_719_0 == 1) v_718_0 <= v_722_0;
      if (v_726_0 == 1) v_725_0 <= v_729_0;
      if (v_733_0 == 1) v_732_0 <= v_736_0;
      if (v_740_0 == 1) v_739_0 <= v_743_0;
      if (v_747_0 == 1) v_746_0 <= v_750_0;
      if (v_754_0 == 1) v_753_0 <= v_757_0;
      if (v_761_0 == 1) v_760_0 <= v_764_0;
      if (v_768_0 == 1) v_767_0 <= v_771_0;
      if (v_775_0 == 1) v_774_0 <= v_778_0;
      if (v_782_0 == 1) v_781_0 <= v_785_0;
      if (v_789_0 == 1) v_788_0 <= v_792_0;
      if (v_796_0 == 1) v_795_0 <= v_799_0;
      if (v_803_0 == 1) v_802_0 <= v_806_0;
      if (v_810_0 == 1) v_809_0 <= v_813_0;
      if (v_817_0 == 1) v_816_0 <= v_820_0;
      if (v_824_0 == 1) v_823_0 <= v_827_0;
      if (v_831_0 == 1) v_830_0 <= v_834_0;
      if (v_838_0 == 1) v_837_0 <= v_841_0;
      if (v_845_0 == 1) v_844_0 <= v_848_0;
      if (v_852_0 == 1) v_851_0 <= v_855_0;
      if (v_859_0 == 1) v_858_0 <= v_862_0;
      if (v_866_0 == 1) v_865_0 <= v_869_0;
      if (v_873_0 == 1) v_872_0 <= v_876_0;
      if (v_880_0 == 1) v_879_0 <= v_883_0;
      if (v_887_0 == 1) v_886_0 <= v_890_0;
      if (v_894_0 == 1) v_893_0 <= v_897_0;
      if (v_901_0 == 1) v_900_0 <= v_904_0;
      if (v_908_0 == 1) v_907_0 <= v_911_0;
      if (v_915_0 == 1) v_914_0 <= v_918_0;
      if (v_922_0 == 1) v_921_0 <= v_925_0;
      if (v_929_0 == 1) v_928_0 <= v_932_0;
      if (v_936_0 == 1) v_935_0 <= v_939_0;
      if (v_943_0 == 1) v_942_0 <= v_946_0;
      if (v_950_0 == 1) v_949_0 <= v_953_0;
      if (v_957_0 == 1) v_956_0 <= v_960_0;
      if (v_964_0 == 1) v_963_0 <= v_967_0;
      if (v_971_0 == 1) v_970_0 <= v_974_0;
      if (v_978_0 == 1) v_977_0 <= v_981_0;
      if (v_985_0 == 1) v_984_0 <= v_988_0;
      if (v_992_0 == 1) v_991_0 <= v_995_0;
      if (v_999_0 == 1) v_998_0 <= v_1002_0;
      if (v_1006_0 == 1) v_1005_0 <= v_1009_0;
      if (v_1013_0 == 1) v_1012_0 <= v_1016_0;
      if (v_1020_0 == 1) v_1019_0 <= v_1023_0;
      if (v_1027_0 == 1) v_1026_0 <= v_1030_0;
      if (v_1034_0 == 1) v_1033_0 <= v_1037_0;
      if (v_1041_0 == 1) v_1040_0 <= v_1044_0;
      if (v_1048_0 == 1) v_1047_0 <= v_1051_0;
      if (v_1055_0 == 1) v_1054_0 <= v_1058_0;
      if (v_1062_0 == 1) v_1061_0 <= v_1065_0;
      if (v_1069_0 == 1) v_1068_0 <= v_1072_0;
      if (v_1076_0 == 1) v_1075_0 <= v_1079_0;
      if (v_1083_0 == 1) v_1082_0 <= v_1086_0;
      if (v_1090_0 == 1) v_1089_0 <= v_1093_0;
      if (v_1097_0 == 1) v_1096_0 <= v_1100_0;
      if (v_1104_0 == 1) v_1103_0 <= v_1107_0;
      if (v_1111_0 == 1) v_1110_0 <= v_1114_0;
      if (v_1118_0 == 1) v_1117_0 <= v_1121_0;
      if (v_1125_0 == 1) v_1124_0 <= v_1128_0;
      if (v_1132_0 == 1) v_1131_0 <= v_1135_0;
      if (v_1139_0 == 1) v_1138_0 <= v_1142_0;
      if (v_1146_0 == 1) v_1145_0 <= v_1149_0;
      if (v_1153_0 == 1) v_1152_0 <= v_1156_0;
      if (v_1160_0 == 1) v_1159_0 <= v_1163_0;
      if (v_1167_0 == 1) v_1166_0 <= v_1170_0;
      if (v_1174_0 == 1) v_1173_0 <= v_1177_0;
      if (v_1181_0 == 1) v_1180_0 <= v_1184_0;
      if (v_1188_0 == 1) v_1187_0 <= v_1191_0;
      if (v_1195_0 == 1) v_1194_0 <= v_1198_0;
      if (v_1202_0 == 1) v_1201_0 <= v_1205_0;
      if (v_1209_0 == 1) v_1208_0 <= v_1212_0;
      if (v_1216_0 == 1) v_1215_0 <= v_1219_0;
      if (v_1223_0 == 1) v_1222_0 <= v_1226_0;
      if (v_1230_0 == 1) v_1229_0 <= v_1233_0;
      if (v_1237_0 == 1) v_1236_0 <= v_1240_0;
      if (v_1244_0 == 1) v_1243_0 <= v_1247_0;
      if (v_1251_0 == 1) v_1250_0 <= v_1254_0;
      if (v_1258_0 == 1) v_1257_0 <= v_1261_0;
      if (v_1265_0 == 1) v_1264_0 <= v_1268_0;
      if (v_1272_0 == 1) v_1271_0 <= v_1275_0;
      if (v_1279_0 == 1) v_1278_0 <= v_1282_0;
      if (v_1286_0 == 1) v_1285_0 <= v_1289_0;
      if (v_1293_0 == 1) v_1292_0 <= v_1296_0;
      if (v_1300_0 == 1) v_1299_0 <= v_1303_0;
      if (v_1307_0 == 1) v_1306_0 <= v_1310_0;
      if (v_1314_0 == 1) v_1313_0 <= v_1317_0;
      if (v_1321_0 == 1) v_1320_0 <= v_1324_0;
      if (v_1328_0 == 1) v_1327_0 <= v_1331_0;
      if (v_1335_0 == 1) v_1334_0 <= v_1338_0;
      if (v_1342_0 == 1) v_1341_0 <= v_1345_0;
      if (v_1349_0 == 1) v_1348_0 <= v_1352_0;
      if (v_1356_0 == 1) v_1355_0 <= v_1359_0;
      if (v_1363_0 == 1) v_1362_0 <= v_1366_0;
      if (v_1370_0 == 1) v_1369_0 <= v_1373_0;
      if (v_1377_0 == 1) v_1376_0 <= v_1380_0;
      if (v_1384_0 == 1) v_1383_0 <= v_1387_0;
      if (v_1391_0 == 1) v_1390_0 <= v_1394_0;
      if (v_1398_0 == 1) v_1397_0 <= v_1401_0;
      if (v_1405_0 == 1) v_1404_0 <= v_1408_0;
      if (v_1412_0 == 1) v_1411_0 <= v_1415_0;
      if (v_1419_0 == 1) v_1418_0 <= v_1422_0;
      if (v_1426_0 == 1) v_1425_0 <= v_1429_0;
      if (v_1433_0 == 1) v_1432_0 <= v_1436_0;
      if (v_1440_0 == 1) v_1439_0 <= v_1443_0;
      if (v_1447_0 == 1) v_1446_0 <= v_1450_0;
      if (v_1454_0 == 1) v_1453_0 <= v_1457_0;
      if (v_1461_0 == 1) v_1460_0 <= v_1464_0;
      if (v_1468_0 == 1) v_1467_0 <= v_1471_0;
      if (v_1475_0 == 1) v_1474_0 <= v_1478_0;
      if (v_1482_0 == 1) v_1481_0 <= v_1485_0;
      if (v_1489_0 == 1) v_1488_0 <= v_1492_0;
      if (v_1496_0 == 1) v_1495_0 <= v_1499_0;
      if (v_1503_0 == 1) v_1502_0 <= v_1506_0;
      if (v_1510_0 == 1) v_1509_0 <= v_1513_0;
      if (v_1517_0 == 1) v_1516_0 <= v_1520_0;
      if (v_1524_0 == 1) v_1523_0 <= v_1527_0;
      if (v_1531_0 == 1) v_1530_0 <= v_1534_0;
      if (v_1538_0 == 1) v_1537_0 <= v_1541_0;
      if (v_1545_0 == 1) v_1544_0 <= v_1548_0;
      if (v_1552_0 == 1) v_1551_0 <= v_1555_0;
      if (v_1559_0 == 1) v_1558_0 <= v_1562_0;
      if (v_1566_0 == 1) v_1565_0 <= v_1569_0;
      if (v_1573_0 == 1) v_1572_0 <= v_1576_0;
      if (v_1580_0 == 1) v_1579_0 <= v_1583_0;
      if (v_1587_0 == 1) v_1586_0 <= v_1590_0;
      if (v_1594_0 == 1) v_1593_0 <= v_1597_0;
      if (v_1601_0 == 1) v_1600_0 <= v_1604_0;
      if (v_1608_0 == 1) v_1607_0 <= v_1611_0;
      if (v_1615_0 == 1) v_1614_0 <= v_1618_0;
      if (v_1622_0 == 1) v_1621_0 <= v_1625_0;
      if (v_1629_0 == 1) v_1628_0 <= v_1632_0;
      if (v_1636_0 == 1) v_1635_0 <= v_1639_0;
      if (v_1643_0 == 1) v_1642_0 <= v_1646_0;
      if (v_1650_0 == 1) v_1649_0 <= v_1653_0;
      if (v_1657_0 == 1) v_1656_0 <= v_1660_0;
      if (v_1664_0 == 1) v_1663_0 <= v_1667_0;
      if (v_1671_0 == 1) v_1670_0 <= v_1674_0;
      if (v_1678_0 == 1) v_1677_0 <= v_1681_0;
      if (v_1685_0 == 1) v_1684_0 <= v_1688_0;
      if (v_1692_0 == 1) v_1691_0 <= v_1695_0;
      if (v_1699_0 == 1) v_1698_0 <= v_1702_0;
      if (v_1706_0 == 1) v_1705_0 <= v_1709_0;
      if (v_1713_0 == 1) v_1712_0 <= v_1716_0;
      if (v_1720_0 == 1) v_1719_0 <= v_1723_0;
      if (v_1727_0 == 1) v_1726_0 <= v_1730_0;
      if (v_1734_0 == 1) v_1733_0 <= v_1737_0;
      if (v_1741_0 == 1) v_1740_0 <= v_1744_0;
      if (v_1748_0 == 1) v_1747_0 <= v_1751_0;
      if (v_1755_0 == 1) v_1754_0 <= v_1758_0;
      if (v_1762_0 == 1) v_1761_0 <= v_1765_0;
      if (v_1769_0 == 1) v_1768_0 <= v_1772_0;
      if (v_1776_0 == 1) v_1775_0 <= v_1779_0;
      if (v_1783_0 == 1) v_1782_0 <= v_1786_0;
      if (v_1790_0 == 1) v_1789_0 <= v_1793_0;
      if (v_1797_0 == 1) v_1796_0 <= v_1800_0;
      if (v_1804_0 == 1) v_1803_0 <= v_1807_0;
      if (v_1811_0 == 1) v_1810_0 <= v_1814_0;
      if (v_1818_0 == 1) v_1817_0 <= v_1821_0;
      if (v_1825_0 == 1) v_1824_0 <= v_1828_0;
      if (v_1832_0 == 1) v_1831_0 <= v_1835_0;
      if (v_1839_0 == 1) v_1838_0 <= v_1842_0;
      if (v_1846_0 == 1) v_1845_0 <= v_1849_0;
      if (v_1853_0 == 1) v_1852_0 <= v_1856_0;
      if (v_1860_0 == 1) v_1859_0 <= v_1863_0;
      if (v_1867_0 == 1) v_1866_0 <= v_1870_0;
      if (v_1874_0 == 1) v_1873_0 <= v_1877_0;
      if (v_1881_0 == 1) v_1880_0 <= v_1884_0;
      if (v_1888_0 == 1) v_1887_0 <= v_1891_0;
      if (v_1895_0 == 1) v_1894_0 <= v_1898_0;
      if (v_1902_0 == 1) v_1901_0 <= v_1905_0;
      if (v_1909_0 == 1) v_1908_0 <= v_1912_0;
      if (v_1916_0 == 1) v_1915_0 <= v_1919_0;
      if (v_1923_0 == 1) v_1922_0 <= v_1926_0;
      if (v_1930_0 == 1) v_1929_0 <= v_1933_0;
      if (v_1937_0 == 1) v_1936_0 <= v_1940_0;
      if (v_1944_0 == 1) v_1943_0 <= v_1947_0;
      if (v_1951_0 == 1) v_1950_0 <= v_1954_0;
      if (v_1958_0 == 1) v_1957_0 <= v_1961_0;
      if (v_1965_0 == 1) v_1964_0 <= v_1968_0;
      if (v_1972_0 == 1) v_1971_0 <= v_1975_0;
      if (v_1979_0 == 1) v_1978_0 <= v_1982_0;
      if (v_1986_0 == 1) v_1985_0 <= v_1989_0;
      if (v_1993_0 == 1) v_1992_0 <= v_1996_0;
      if (v_2000_0 == 1) v_1999_0 <= v_2003_0;
      if (v_2007_0 == 1) v_2006_0 <= v_2010_0;
      if (v_2014_0 == 1) v_2013_0 <= v_2017_0;
      if (v_2021_0 == 1) v_2020_0 <= v_2024_0;
      if (v_2028_0 == 1) v_2027_0 <= v_2031_0;
      if (v_2035_0 == 1) v_2034_0 <= v_2038_0;
      if (v_2042_0 == 1) v_2041_0 <= v_2045_0;
      if (v_2049_0 == 1) v_2048_0 <= v_2052_0;
      if (v_2056_0 == 1) v_2055_0 <= v_2059_0;
      if (v_2063_0 == 1) v_2062_0 <= v_2066_0;
      if (v_2070_0 == 1) v_2069_0 <= v_2073_0;
      if (v_2077_0 == 1) v_2076_0 <= v_2080_0;
      if (v_2084_0 == 1) v_2083_0 <= v_2087_0;
      if (v_2091_0 == 1) v_2090_0 <= v_2094_0;
      if (v_2098_0 == 1) v_2097_0 <= v_2101_0;
      if (v_2105_0 == 1) v_2104_0 <= v_2108_0;
      if (v_2112_0 == 1) v_2111_0 <= v_2115_0;
      if (v_2119_0 == 1) v_2118_0 <= v_2122_0;
      if (v_2126_0 == 1) v_2125_0 <= v_2129_0;
      if (v_2133_0 == 1) v_2132_0 <= v_2136_0;
      if (v_2140_0 == 1) v_2139_0 <= v_2143_0;
      if (v_2147_0 == 1) v_2146_0 <= v_2150_0;
      if (v_2154_0 == 1) v_2153_0 <= v_2157_0;
      if (v_2161_0 == 1) v_2160_0 <= v_2164_0;
      if (v_2168_0 == 1) v_2167_0 <= v_2171_0;
      if (v_2175_0 == 1) v_2174_0 <= v_2178_0;
      if (v_2182_0 == 1) v_2181_0 <= v_2185_0;
      if (v_2189_0 == 1) v_2188_0 <= v_2192_0;
      if (v_2196_0 == 1) v_2195_0 <= v_2199_0;
      if (v_2203_0 == 1) v_2202_0 <= v_2206_0;
      if (v_2210_0 == 1) v_2209_0 <= v_2213_0;
      if (v_2217_0 == 1) v_2216_0 <= v_2220_0;
      if (v_2224_0 == 1) v_2223_0 <= v_2227_0;
      if (v_2231_0 == 1) v_2230_0 <= v_2234_0;
      if (v_2238_0 == 1) v_2237_0 <= v_2241_0;
      if (v_2245_0 == 1) v_2244_0 <= v_2248_0;
      if (v_2252_0 == 1) v_2251_0 <= v_2255_0;
      if (v_2259_0 == 1) v_2258_0 <= v_2262_0;
      if (v_2266_0 == 1) v_2265_0 <= v_2269_0;
      if (v_2273_0 == 1) v_2272_0 <= v_2276_0;
      if (v_2280_0 == 1) v_2279_0 <= v_2283_0;
      if (v_2287_0 == 1) v_2286_0 <= v_2290_0;
      if (v_2294_0 == 1) v_2293_0 <= v_2297_0;
      if (v_2301_0 == 1) v_2300_0 <= v_2304_0;
      if (v_2308_0 == 1) v_2307_0 <= v_2311_0;
      if (v_2315_0 == 1) v_2314_0 <= v_2318_0;
      if (v_2322_0 == 1) v_2321_0 <= v_2325_0;
      if (v_2329_0 == 1) v_2328_0 <= v_2332_0;
      if (v_2336_0 == 1) v_2335_0 <= v_2339_0;
      if (v_2343_0 == 1) v_2342_0 <= v_2346_0;
      if (v_2350_0 == 1) v_2349_0 <= v_2353_0;
      if (v_2357_0 == 1) v_2356_0 <= v_2360_0;
      if (v_2364_0 == 1) v_2363_0 <= v_2367_0;
      if (v_2371_0 == 1) v_2370_0 <= v_2374_0;
      if (v_2378_0 == 1) v_2377_0 <= v_2381_0;
      if (v_2385_0 == 1) v_2384_0 <= v_2388_0;
      if (v_2392_0 == 1) v_2391_0 <= v_2395_0;
      if (v_2399_0 == 1) v_2398_0 <= v_2402_0;
      if (v_2406_0 == 1) v_2405_0 <= v_2409_0;
      if (v_2413_0 == 1) v_2412_0 <= v_2416_0;
      if (v_2420_0 == 1) v_2419_0 <= v_2423_0;
      if (v_2427_0 == 1) v_2426_0 <= v_2430_0;
      if (v_2434_0 == 1) v_2433_0 <= v_2437_0;
      if (v_2441_0 == 1) v_2440_0 <= v_2444_0;
      if (v_2448_0 == 1) v_2447_0 <= v_2451_0;
      if (v_2455_0 == 1) v_2454_0 <= v_2458_0;
      if (v_2462_0 == 1) v_2461_0 <= v_2465_0;
      if (v_2469_0 == 1) v_2468_0 <= v_2472_0;
      if (v_2476_0 == 1) v_2475_0 <= v_2479_0;
      if (v_2483_0 == 1) v_2482_0 <= v_2486_0;
      if (v_2490_0 == 1) v_2489_0 <= v_2493_0;
      if (v_2497_0 == 1) v_2496_0 <= v_2500_0;
      if (v_2504_0 == 1) v_2503_0 <= v_2507_0;
      if (v_2511_0 == 1) v_2510_0 <= v_2514_0;
      if (v_2518_0 == 1) v_2517_0 <= v_2521_0;
      if (v_2525_0 == 1) v_2524_0 <= v_2528_0;
      if (v_2532_0 == 1) v_2531_0 <= v_2535_0;
      if (v_2539_0 == 1) v_2538_0 <= v_2542_0;
      if (v_2546_0 == 1) v_2545_0 <= v_2549_0;
      if (v_2553_0 == 1) v_2552_0 <= v_2556_0;
      if (v_2560_0 == 1) v_2559_0 <= v_2563_0;
      if (v_2567_0 == 1) v_2566_0 <= v_2570_0;
      if (v_2574_0 == 1) v_2573_0 <= v_2577_0;
      if (v_2581_0 == 1) v_2580_0 <= v_2584_0;
      if (v_2588_0 == 1) v_2587_0 <= v_2591_0;
      if (v_2595_0 == 1) v_2594_0 <= v_2598_0;
      if (v_2602_0 == 1) v_2601_0 <= v_2605_0;
      if (v_2609_0 == 1) v_2608_0 <= v_2612_0;
      if (v_2616_0 == 1) v_2615_0 <= v_2619_0;
      if (v_2623_0 == 1) v_2622_0 <= v_2626_0;
      if (v_2630_0 == 1) v_2629_0 <= v_2633_0;
      if (v_2637_0 == 1) v_2636_0 <= v_2640_0;
      if (v_2644_0 == 1) v_2643_0 <= v_2647_0;
      if (v_2651_0 == 1) v_2650_0 <= v_2654_0;
      if (v_2658_0 == 1) v_2657_0 <= v_2661_0;
      if (v_2665_0 == 1) v_2664_0 <= v_2668_0;
      if (v_2672_0 == 1) v_2671_0 <= v_2675_0;
      if (v_2679_0 == 1) v_2678_0 <= v_2682_0;
      if (v_2686_0 == 1) v_2685_0 <= v_2689_0;
      if (v_2693_0 == 1) v_2692_0 <= v_2696_0;
      if (v_2700_0 == 1) v_2699_0 <= v_2703_0;
      if (v_2707_0 == 1) v_2706_0 <= v_2710_0;
      if (v_2714_0 == 1) v_2713_0 <= v_2717_0;
      if (v_2721_0 == 1) v_2720_0 <= v_2724_0;
      if (v_2728_0 == 1) v_2727_0 <= v_2731_0;
      if (v_2735_0 == 1) v_2734_0 <= v_2738_0;
      if (v_2742_0 == 1) v_2741_0 <= v_2745_0;
      if (v_2749_0 == 1) v_2748_0 <= v_2752_0;
      if (v_2756_0 == 1) v_2755_0 <= v_2759_0;
      if (v_2763_0 == 1) v_2762_0 <= v_2766_0;
      if (v_2770_0 == 1) v_2769_0 <= v_2773_0;
      if (v_2777_0 == 1) v_2776_0 <= v_2780_0;
      if (v_2784_0 == 1) v_2783_0 <= v_2787_0;
      if (v_2791_0 == 1) v_2790_0 <= v_2794_0;
      if (v_2798_0 == 1) v_2797_0 <= v_2801_0;
      if (v_2805_0 == 1) v_2804_0 <= v_2808_0;
      if (v_2812_0 == 1) v_2811_0 <= v_2815_0;
      if (v_2819_0 == 1) v_2818_0 <= v_2822_0;
      if (v_2826_0 == 1) v_2825_0 <= v_2829_0;
      if (v_2833_0 == 1) v_2832_0 <= v_2836_0;
      if (v_2840_0 == 1) v_2839_0 <= v_2843_0;
      if (v_2847_0 == 1) v_2846_0 <= v_2850_0;
      if (v_2854_0 == 1) v_2853_0 <= v_2857_0;
      if (v_2861_0 == 1) v_2860_0 <= v_2864_0;
      if (v_2868_0 == 1) v_2867_0 <= v_2871_0;
      if (v_2875_0 == 1) v_2874_0 <= v_2878_0;
      if (v_2882_0 == 1) v_2881_0 <= v_2885_0;
      if (v_2889_0 == 1) v_2888_0 <= v_2892_0;
      if (v_2896_0 == 1) v_2895_0 <= v_2899_0;
      if (v_2903_0 == 1) v_2902_0 <= v_2906_0;
      if (v_2910_0 == 1) v_2909_0 <= v_2913_0;
      if (v_2917_0 == 1) v_2916_0 <= v_2920_0;
      if (v_2924_0 == 1) v_2923_0 <= v_2927_0;
      if (v_2931_0 == 1) v_2930_0 <= v_2934_0;
      if (v_2938_0 == 1) v_2937_0 <= v_2941_0;
      if (v_2945_0 == 1) v_2944_0 <= v_2948_0;
      if (v_2952_0 == 1) v_2951_0 <= v_2955_0;
      if (v_2959_0 == 1) v_2958_0 <= v_2962_0;
      if (v_2966_0 == 1) v_2965_0 <= v_2969_0;
      if (v_2973_0 == 1) v_2972_0 <= v_2976_0;
      if (v_2980_0 == 1) v_2979_0 <= v_2983_0;
      if (v_2987_0 == 1) v_2986_0 <= v_2990_0;
      if (v_2994_0 == 1) v_2993_0 <= v_2997_0;
      if (v_3001_0 == 1) v_3000_0 <= v_3004_0;
      if (v_3008_0 == 1) v_3007_0 <= v_3011_0;
      if (v_3015_0 == 1) v_3014_0 <= v_3018_0;
      if (v_3022_0 == 1) v_3021_0 <= v_3025_0;
      if (v_3029_0 == 1) v_3028_0 <= v_3032_0;
      if (v_3036_0 == 1) v_3035_0 <= v_3039_0;
      if (v_3043_0 == 1) v_3042_0 <= v_3046_0;
      if (v_3050_0 == 1) v_3049_0 <= v_3053_0;
      if (v_3057_0 == 1) v_3056_0 <= v_3060_0;
      if (v_3064_0 == 1) v_3063_0 <= v_3067_0;
      if (v_3071_0 == 1) v_3070_0 <= v_3074_0;
      if (v_3078_0 == 1) v_3077_0 <= v_3081_0;
      if (v_3085_0 == 1) v_3084_0 <= v_3088_0;
      if (v_3092_0 == 1) v_3091_0 <= v_3095_0;
      if (v_3099_0 == 1) v_3098_0 <= v_3102_0;
      if (v_3106_0 == 1) v_3105_0 <= v_3109_0;
      if (v_3113_0 == 1) v_3112_0 <= v_3116_0;
      if (v_3120_0 == 1) v_3119_0 <= v_3123_0;
      if (v_3127_0 == 1) v_3126_0 <= v_3130_0;
      if (v_3134_0 == 1) v_3133_0 <= v_3137_0;
      if (v_3141_0 == 1) v_3140_0 <= v_3144_0;
      if (v_3148_0 == 1) v_3147_0 <= v_3151_0;
      if (v_3155_0 == 1) v_3154_0 <= v_3158_0;
      if (v_3162_0 == 1) v_3161_0 <= v_3165_0;
      if (v_3169_0 == 1) v_3168_0 <= v_3172_0;
      if (v_3176_0 == 1) v_3175_0 <= v_3179_0;
      if (v_3183_0 == 1) v_3182_0 <= v_3186_0;
      if (v_3190_0 == 1) v_3189_0 <= v_3193_0;
      if (v_3197_0 == 1) v_3196_0 <= v_3200_0;
      if (v_3204_0 == 1) v_3203_0 <= v_3207_0;
      if (v_3211_0 == 1) v_3210_0 <= v_3214_0;
      if (v_3218_0 == 1) v_3217_0 <= v_3221_0;
      if (v_3225_0 == 1) v_3224_0 <= v_3228_0;
      if (v_3232_0 == 1) v_3231_0 <= v_3235_0;
      if (v_3239_0 == 1) v_3238_0 <= v_3242_0;
      if (v_3246_0 == 1) v_3245_0 <= v_3249_0;
      if (v_3253_0 == 1) v_3252_0 <= v_3256_0;
      if (v_3260_0 == 1) v_3259_0 <= v_3263_0;
      if (v_3267_0 == 1) v_3266_0 <= v_3270_0;
      if (v_3274_0 == 1) v_3273_0 <= v_3277_0;
      if (v_3281_0 == 1) v_3280_0 <= v_3284_0;
      if (v_3288_0 == 1) v_3287_0 <= v_3291_0;
      if (v_3295_0 == 1) v_3294_0 <= v_3298_0;
      if (v_3302_0 == 1) v_3301_0 <= v_3305_0;
      if (v_3309_0 == 1) v_3308_0 <= v_3312_0;
      if (v_3316_0 == 1) v_3315_0 <= v_3319_0;
      if (v_3323_0 == 1) v_3322_0 <= v_3326_0;
      if (v_3330_0 == 1) v_3329_0 <= v_3333_0;
      if (v_3337_0 == 1) v_3336_0 <= v_3340_0;
      if (v_3344_0 == 1) v_3343_0 <= v_3347_0;
      if (v_3351_0 == 1) v_3350_0 <= v_3354_0;
      if (v_3358_0 == 1) v_3357_0 <= v_3361_0;
      if (v_3365_0 == 1) v_3364_0 <= v_3368_0;
      if (v_3372_0 == 1) v_3371_0 <= v_3375_0;
      if (v_3379_0 == 1) v_3378_0 <= v_3382_0;
      if (v_3386_0 == 1) v_3385_0 <= v_3389_0;
      if (v_3393_0 == 1) v_3392_0 <= v_3396_0;
      if (v_3400_0 == 1) v_3399_0 <= v_3403_0;
      if (v_3407_0 == 1) v_3406_0 <= v_3410_0;
      if (v_3414_0 == 1) v_3413_0 <= v_3417_0;
      if (v_3421_0 == 1) v_3420_0 <= v_3424_0;
      if (v_3428_0 == 1) v_3427_0 <= v_3431_0;
      if (v_3435_0 == 1) v_3434_0 <= v_3438_0;
      if (v_3442_0 == 1) v_3441_0 <= v_3445_0;
      if (v_3449_0 == 1) v_3448_0 <= v_3452_0;
      if (v_3456_0 == 1) v_3455_0 <= v_3459_0;
      if (v_3463_0 == 1) v_3462_0 <= v_3466_0;
      if (v_3470_0 == 1) v_3469_0 <= v_3473_0;
      if (v_3477_0 == 1) v_3476_0 <= v_3480_0;
      if (v_3484_0 == 1) v_3483_0 <= v_3487_0;
      if (v_3491_0 == 1) v_3490_0 <= v_3494_0;
      if (v_3498_0 == 1) v_3497_0 <= v_3501_0;
      if (v_3505_0 == 1) v_3504_0 <= v_3508_0;
      if (v_3512_0 == 1) v_3511_0 <= v_3515_0;
      if (v_3519_0 == 1) v_3518_0 <= v_3522_0;
      if (v_3526_0 == 1) v_3525_0 <= v_3529_0;
      if (v_3533_0 == 1) v_3532_0 <= v_3536_0;
      if (v_3540_0 == 1) v_3539_0 <= v_3543_0;
      if (v_3547_0 == 1) v_3546_0 <= v_3550_0;
      if (v_3554_0 == 1) v_3553_0 <= v_3557_0;
      if (v_3561_0 == 1) v_3560_0 <= v_3564_0;
      if (v_3568_0 == 1) v_3567_0 <= v_3571_0;
      if (v_3575_0 == 1) v_3574_0 <= v_3578_0;
      if (v_3582_0 == 1) v_3581_0 <= v_3585_0;
      if (v_3589_0 == 1) v_3588_0 <= v_3592_0;
      if (v_3596_0 == 1) v_3595_0 <= v_3599_0;
      if (v_3603_0 == 1) v_3602_0 <= v_3606_0;
      if (v_3610_0 == 1) v_3609_0 <= v_3613_0;
      if (v_3617_0 == 1) v_3616_0 <= v_3620_0;
      if (v_3624_0 == 1) v_3623_0 <= v_3627_0;
      if (v_3631_0 == 1) v_3630_0 <= v_3634_0;
      if (v_3638_0 == 1) v_3637_0 <= v_3641_0;
      if (v_3645_0 == 1) v_3644_0 <= v_3648_0;
      if (v_3652_0 == 1) v_3651_0 <= v_3655_0;
      if (v_3659_0 == 1) v_3658_0 <= v_3662_0;
      if (v_3666_0 == 1) v_3665_0 <= v_3669_0;
      if (v_3673_0 == 1) v_3672_0 <= v_3676_0;
      if (v_3680_0 == 1) v_3679_0 <= v_3683_0;
      if (v_3687_0 == 1) v_3686_0 <= v_3690_0;
      if (v_3694_0 == 1) v_3693_0 <= v_3697_0;
      if (v_3701_0 == 1) v_3700_0 <= v_3704_0;
      if (v_3708_0 == 1) v_3707_0 <= v_3711_0;
      if (v_3715_0 == 1) v_3714_0 <= v_3718_0;
      if (v_3722_0 == 1) v_3721_0 <= v_3725_0;
      if (v_3729_0 == 1) v_3728_0 <= v_3732_0;
      if (v_3736_0 == 1) v_3735_0 <= v_3739_0;
      if (v_3743_0 == 1) v_3742_0 <= v_3746_0;
      if (v_3750_0 == 1) v_3749_0 <= v_3753_0;
      if (v_3757_0 == 1) v_3756_0 <= v_3760_0;
      if (v_3764_0 == 1) v_3763_0 <= v_3767_0;
      if (v_3771_0 == 1) v_3770_0 <= v_3774_0;
      if (v_3778_0 == 1) v_3777_0 <= v_3781_0;
      if (v_3785_0 == 1) v_3784_0 <= v_3788_0;
      if (v_3792_0 == 1) v_3791_0 <= v_3795_0;
      if (v_3799_0 == 1) v_3798_0 <= v_3802_0;
      if (v_3806_0 == 1) v_3805_0 <= v_3809_0;
      if (v_3813_0 == 1) v_3812_0 <= v_3816_0;
      if (v_3820_0 == 1) v_3819_0 <= v_3823_0;
      if (v_3827_0 == 1) v_3826_0 <= v_3830_0;
      if (v_3834_0 == 1) v_3833_0 <= v_3837_0;
      if (v_3841_0 == 1) v_3840_0 <= v_3844_0;
      if (v_3848_0 == 1) v_3847_0 <= v_3851_0;
      if (v_3855_0 == 1) v_3854_0 <= v_3858_0;
      if (v_3862_0 == 1) v_3861_0 <= v_3865_0;
      if (v_3869_0 == 1) v_3868_0 <= v_3872_0;
      if (v_3876_0 == 1) v_3875_0 <= v_3879_0;
      if (v_3883_0 == 1) v_3882_0 <= v_3886_0;
      if (v_3890_0 == 1) v_3889_0 <= v_3893_0;
      if (v_3897_0 == 1) v_3896_0 <= v_3900_0;
      if (v_3904_0 == 1) v_3903_0 <= v_3907_0;
      if (v_3911_0 == 1) v_3910_0 <= v_3914_0;
      if (v_3918_0 == 1) v_3917_0 <= v_3921_0;
      if (v_3925_0 == 1) v_3924_0 <= v_3928_0;
      if (v_3932_0 == 1) v_3931_0 <= v_3935_0;
      if (v_3939_0 == 1) v_3938_0 <= v_3942_0;
      if (v_3946_0 == 1) v_3945_0 <= v_3949_0;
      if (v_3953_0 == 1) v_3952_0 <= v_3956_0;
      if (v_3960_0 == 1) v_3959_0 <= v_3963_0;
      if (v_3967_0 == 1) v_3966_0 <= v_3970_0;
      if (v_3974_0 == 1) v_3973_0 <= v_3977_0;
      if (v_3981_0 == 1) v_3980_0 <= v_3984_0;
      if (v_3988_0 == 1) v_3987_0 <= v_3991_0;
      if (v_3995_0 == 1) v_3994_0 <= v_3998_0;
      if (v_4002_0 == 1) v_4001_0 <= v_4005_0;
      if (v_4009_0 == 1) v_4008_0 <= v_4012_0;
      if (v_4016_0 == 1) v_4015_0 <= v_4019_0;
      if (v_4023_0 == 1) v_4022_0 <= v_4026_0;
      if (v_4030_0 == 1) v_4029_0 <= v_4033_0;
      if (v_4037_0 == 1) v_4036_0 <= v_4040_0;
      if (v_4044_0 == 1) v_4043_0 <= v_4047_0;
      if (v_4051_0 == 1) v_4050_0 <= v_4054_0;
      if (v_4058_0 == 1) v_4057_0 <= v_4061_0;
      if (v_4065_0 == 1) v_4064_0 <= v_4068_0;
      if (v_4072_0 == 1) v_4071_0 <= v_4075_0;
      if (v_4079_0 == 1) v_4078_0 <= v_4082_0;
      if (v_4086_0 == 1) v_4085_0 <= v_4089_0;
      if (v_4093_0 == 1) v_4092_0 <= v_4096_0;
      if (v_4100_0 == 1) v_4099_0 <= v_4103_0;
      if (v_4107_0 == 1) v_4106_0 <= v_4110_0;
      if (v_4114_0 == 1) v_4113_0 <= v_4117_0;
      if (v_4121_0 == 1) v_4120_0 <= v_4124_0;
      if (v_4128_0 == 1) v_4127_0 <= v_4131_0;
      if (v_4135_0 == 1) v_4134_0 <= v_4138_0;
      if (v_4142_0 == 1) v_4141_0 <= v_4145_0;
      if (v_4149_0 == 1) v_4148_0 <= v_4152_0;
      if (v_4156_0 == 1) v_4155_0 <= v_4159_0;
      if (v_4163_0 == 1) v_4162_0 <= v_4166_0;
      if (v_4170_0 == 1) v_4169_0 <= v_4173_0;
      if (v_4177_0 == 1) v_4176_0 <= v_4180_0;
      if (v_4184_0 == 1) v_4183_0 <= v_4187_0;
      if (v_4191_0 == 1) v_4190_0 <= v_4194_0;
      if (v_4198_0 == 1) v_4197_0 <= v_4201_0;
      if (v_4205_0 == 1) v_4204_0 <= v_4208_0;
      if (v_4212_0 == 1) v_4211_0 <= v_4215_0;
      if (v_4219_0 == 1) v_4218_0 <= v_4222_0;
      if (v_4226_0 == 1) v_4225_0 <= v_4229_0;
      if (v_4233_0 == 1) v_4232_0 <= v_4236_0;
      if (v_4240_0 == 1) v_4239_0 <= v_4243_0;
      if (v_4247_0 == 1) v_4246_0 <= v_4250_0;
      if (v_4254_0 == 1) v_4253_0 <= v_4257_0;
      if (v_4261_0 == 1) v_4260_0 <= v_4264_0;
      if (v_4268_0 == 1) v_4267_0 <= v_4271_0;
      if (v_4275_0 == 1) v_4274_0 <= v_4278_0;
      if (v_4282_0 == 1) v_4281_0 <= v_4285_0;
      if (v_4289_0 == 1) v_4288_0 <= v_4292_0;
      if (v_4296_0 == 1) v_4295_0 <= v_4299_0;
      if (v_4303_0 == 1) v_4302_0 <= v_4306_0;
      if (v_4310_0 == 1) v_4309_0 <= v_4313_0;
      if (v_4317_0 == 1) v_4316_0 <= v_4320_0;
      if (v_4324_0 == 1) v_4323_0 <= v_4327_0;
      if (v_4331_0 == 1) v_4330_0 <= v_4334_0;
      if (v_4338_0 == 1) v_4337_0 <= v_4341_0;
      if (v_4345_0 == 1) v_4344_0 <= v_4348_0;
      if (v_4352_0 == 1) v_4351_0 <= v_4355_0;
      if (v_4359_0 == 1) v_4358_0 <= v_4362_0;
      if (v_4366_0 == 1) v_4365_0 <= v_4369_0;
      if (v_4373_0 == 1) v_4372_0 <= v_4376_0;
      if (v_4380_0 == 1) v_4379_0 <= v_4383_0;
      if (v_4387_0 == 1) v_4386_0 <= v_4390_0;
      if (v_4394_0 == 1) v_4393_0 <= v_4397_0;
      if (v_4401_0 == 1) v_4400_0 <= v_4404_0;
      if (v_4408_0 == 1) v_4407_0 <= v_4411_0;
      if (v_4415_0 == 1) v_4414_0 <= v_4418_0;
      if (v_4422_0 == 1) v_4421_0 <= v_4425_0;
      if (v_4429_0 == 1) v_4428_0 <= v_4432_0;
      if (v_4436_0 == 1) v_4435_0 <= v_4439_0;
      if (v_4443_0 == 1) v_4442_0 <= v_4446_0;
      if (v_4450_0 == 1) v_4449_0 <= v_4453_0;
      if (v_4457_0 == 1) v_4456_0 <= v_4460_0;
      if (v_4464_0 == 1) v_4463_0 <= v_4467_0;
      if (v_4471_0 == 1) v_4470_0 <= v_4474_0;
      if (v_4478_0 == 1) v_4477_0 <= v_4481_0;
      if (v_4485_0 == 1) v_4484_0 <= v_4488_0;
      if (v_4492_0 == 1) v_4491_0 <= v_4495_0;
      if (v_4499_0 == 1) v_4498_0 <= v_4502_0;
      if (v_4506_0 == 1) v_4505_0 <= v_4509_0;
      if (v_4513_0 == 1) v_4512_0 <= v_4516_0;
      if (v_4520_0 == 1) v_4519_0 <= v_4523_0;
      if (v_4527_0 == 1) v_4526_0 <= v_4530_0;
      if (v_4534_0 == 1) v_4533_0 <= v_4537_0;
      if (v_4541_0 == 1) v_4540_0 <= v_4544_0;
      if (v_4548_0 == 1) v_4547_0 <= v_4551_0;
      if (v_4555_0 == 1) v_4554_0 <= v_4558_0;
      if (v_4562_0 == 1) v_4561_0 <= v_4565_0;
      if (v_4569_0 == 1) v_4568_0 <= v_4572_0;
      if (v_4576_0 == 1) v_4575_0 <= v_4579_0;
      if (v_4583_0 == 1) v_4582_0 <= v_4586_0;
      if (v_4590_0 == 1) v_4589_0 <= v_4593_0;
      if (v_4597_0 == 1) v_4596_0 <= v_4600_0;
      if (v_4604_0 == 1) v_4603_0 <= v_4607_0;
      if (v_4611_0 == 1) v_4610_0 <= v_4614_0;
      if (v_4618_0 == 1) v_4617_0 <= v_4621_0;
      if (v_4625_0 == 1) v_4624_0 <= v_4628_0;
      if (v_4632_0 == 1) v_4631_0 <= v_4635_0;
      if (v_4639_0 == 1) v_4638_0 <= v_4642_0;
      if (v_4646_0 == 1) v_4645_0 <= v_4649_0;
      if (v_4653_0 == 1) v_4652_0 <= v_4656_0;
      if (v_4660_0 == 1) v_4659_0 <= v_4663_0;
      if (v_4667_0 == 1) v_4666_0 <= v_4670_0;
      if (v_4674_0 == 1) v_4673_0 <= v_4677_0;
      if (v_4681_0 == 1) v_4680_0 <= v_4684_0;
      if (v_4688_0 == 1) v_4687_0 <= v_4691_0;
      if (v_4695_0 == 1) v_4694_0 <= v_4698_0;
      if (v_4702_0 == 1) v_4701_0 <= v_4705_0;
      if (v_4709_0 == 1) v_4708_0 <= v_4712_0;
      if (v_4716_0 == 1) v_4715_0 <= v_4719_0;
      if (v_4723_0 == 1) v_4722_0 <= v_4726_0;
      if (v_4730_0 == 1) v_4729_0 <= v_4733_0;
      if (v_4737_0 == 1) v_4736_0 <= v_4740_0;
      if (v_4744_0 == 1) v_4743_0 <= v_4747_0;
      if (v_4751_0 == 1) v_4750_0 <= v_4754_0;
      if (v_4758_0 == 1) v_4757_0 <= v_4761_0;
      if (v_4765_0 == 1) v_4764_0 <= v_4768_0;
      if (v_4772_0 == 1) v_4771_0 <= v_4775_0;
      if (v_4779_0 == 1) v_4778_0 <= v_4782_0;
      if (v_4786_0 == 1) v_4785_0 <= v_4789_0;
      if (v_4793_0 == 1) v_4792_0 <= v_4796_0;
      if (v_4800_0 == 1) v_4799_0 <= v_4803_0;
      if (v_4807_0 == 1) v_4806_0 <= v_4810_0;
      if (v_4814_0 == 1) v_4813_0 <= v_4817_0;
      if (v_4821_0 == 1) v_4820_0 <= v_4824_0;
      if (v_4828_0 == 1) v_4827_0 <= v_4831_0;
      if (v_4835_0 == 1) v_4834_0 <= v_4838_0;
      if (v_4842_0 == 1) v_4841_0 <= v_4845_0;
      if (v_4849_0 == 1) v_4848_0 <= v_4852_0;
      if (v_4856_0 == 1) v_4855_0 <= v_4859_0;
      if (v_4863_0 == 1) v_4862_0 <= v_4866_0;
      if (v_4870_0 == 1) v_4869_0 <= v_4873_0;
      if (v_4877_0 == 1) v_4876_0 <= v_4880_0;
      if (v_4884_0 == 1) v_4883_0 <= v_4887_0;
      if (v_4891_0 == 1) v_4890_0 <= v_4894_0;
      if (v_4898_0 == 1) v_4897_0 <= v_4901_0;
      if (v_4905_0 == 1) v_4904_0 <= v_4908_0;
      if (v_4912_0 == 1) v_4911_0 <= v_4915_0;
      if (v_4919_0 == 1) v_4918_0 <= v_4922_0;
      if (v_4926_0 == 1) v_4925_0 <= v_4929_0;
      if (v_4933_0 == 1) v_4932_0 <= v_4936_0;
      if (v_4940_0 == 1) v_4939_0 <= v_4943_0;
      if (v_4947_0 == 1) v_4946_0 <= v_4950_0;
      if (v_4954_0 == 1) v_4953_0 <= v_4957_0;
      if (v_4961_0 == 1) v_4960_0 <= v_4964_0;
      if (v_4968_0 == 1) v_4967_0 <= v_4971_0;
      if (v_4975_0 == 1) v_4974_0 <= v_4978_0;
      if (v_4982_0 == 1) v_4981_0 <= v_4985_0;
      if (v_4989_0 == 1) v_4988_0 <= v_4992_0;
      if (v_4996_0 == 1) v_4995_0 <= v_4999_0;
      if (v_5003_0 == 1) v_5002_0 <= v_5006_0;
      if (v_5010_0 == 1) v_5009_0 <= v_5013_0;
      if (v_5017_0 == 1) v_5016_0 <= v_5020_0;
      if (v_5024_0 == 1) v_5023_0 <= v_5027_0;
      if (v_5031_0 == 1) v_5030_0 <= v_5034_0;
      if (v_5038_0 == 1) v_5037_0 <= v_5041_0;
      if (v_5045_0 == 1) v_5044_0 <= v_5048_0;
      if (v_5052_0 == 1) v_5051_0 <= v_5055_0;
      if (v_5059_0 == 1) v_5058_0 <= v_5062_0;
      if (v_5066_0 == 1) v_5065_0 <= v_5069_0;
      if (v_5073_0 == 1) v_5072_0 <= v_5076_0;
      if (v_5080_0 == 1) v_5079_0 <= v_5083_0;
      if (v_5087_0 == 1) v_5086_0 <= v_5090_0;
      if (v_5094_0 == 1) v_5093_0 <= v_5097_0;
      if (v_5101_0 == 1) v_5100_0 <= v_5104_0;
      if (v_5108_0 == 1) v_5107_0 <= v_5111_0;
      if (v_5115_0 == 1) v_5114_0 <= v_5118_0;
      if (v_5122_0 == 1) v_5121_0 <= v_5125_0;
      if (v_5129_0 == 1) v_5128_0 <= v_5132_0;
      if (v_5136_0 == 1) v_5135_0 <= v_5139_0;
      if (v_5143_0 == 1) v_5142_0 <= v_5146_0;
      if (v_5150_0 == 1) v_5149_0 <= v_5153_0;
      if (v_5157_0 == 1) v_5156_0 <= v_5160_0;
      if (v_5164_0 == 1) v_5163_0 <= v_5167_0;
      if (v_5171_0 == 1) v_5170_0 <= v_5174_0;
      if (v_5178_0 == 1) v_5177_0 <= v_5181_0;
      if (v_5185_0 == 1) v_5184_0 <= v_5188_0;
      if (v_5192_0 == 1) v_5191_0 <= v_5195_0;
      if (v_5199_0 == 1) v_5198_0 <= v_5202_0;
      if (v_5206_0 == 1) v_5205_0 <= v_5209_0;
      if (v_5213_0 == 1) v_5212_0 <= v_5216_0;
      if (v_5220_0 == 1) v_5219_0 <= v_5223_0;
      if (v_5227_0 == 1) v_5226_0 <= v_5230_0;
      if (v_5234_0 == 1) v_5233_0 <= v_5237_0;
      if (v_5241_0 == 1) v_5240_0 <= v_5244_0;
      if (v_5248_0 == 1) v_5247_0 <= v_5251_0;
      if (v_5255_0 == 1) v_5254_0 <= v_5258_0;
      if (v_5262_0 == 1) v_5261_0 <= v_5265_0;
      if (v_5269_0 == 1) v_5268_0 <= v_5272_0;
      if (v_5276_0 == 1) v_5275_0 <= v_5279_0;
      if (v_5283_0 == 1) v_5282_0 <= v_5286_0;
      if (v_5290_0 == 1) v_5289_0 <= v_5293_0;
      if (v_5297_0 == 1) v_5296_0 <= v_5300_0;
      if (v_5304_0 == 1) v_5303_0 <= v_5307_0;
      if (v_5311_0 == 1) v_5310_0 <= v_5314_0;
      if (v_5318_0 == 1) v_5317_0 <= v_5321_0;
      if (v_5325_0 == 1) v_5324_0 <= v_5328_0;
      if (v_5332_0 == 1) v_5331_0 <= v_5335_0;
      if (v_5339_0 == 1) v_5338_0 <= v_5342_0;
      if (v_5346_0 == 1) v_5345_0 <= v_5349_0;
      if (v_5353_0 == 1) v_5352_0 <= v_5356_0;
      if (v_5360_0 == 1) v_5359_0 <= v_5363_0;
      if (v_5367_0 == 1) v_5366_0 <= v_5370_0;
      if (v_5374_0 == 1) v_5373_0 <= v_5377_0;
      if (v_5381_0 == 1) v_5380_0 <= v_5384_0;
      if (v_5388_0 == 1) v_5387_0 <= v_5391_0;
      if (v_5395_0 == 1) v_5394_0 <= v_5398_0;
      if (v_5402_0 == 1) v_5401_0 <= v_5405_0;
      if (v_5409_0 == 1) v_5408_0 <= v_5412_0;
      if (v_5416_0 == 1) v_5415_0 <= v_5419_0;
      if (v_5423_0 == 1) v_5422_0 <= v_5426_0;
      if (v_5430_0 == 1) v_5429_0 <= v_5433_0;
      if (v_5437_0 == 1) v_5436_0 <= v_5440_0;
      if (v_5444_0 == 1) v_5443_0 <= v_5447_0;
      if (v_5451_0 == 1) v_5450_0 <= v_5454_0;
      if (v_5458_0 == 1) v_5457_0 <= v_5461_0;
      if (v_5465_0 == 1) v_5464_0 <= v_5468_0;
      if (v_5472_0 == 1) v_5471_0 <= v_5475_0;
      if (v_5479_0 == 1) v_5478_0 <= v_5482_0;
      if (v_5486_0 == 1) v_5485_0 <= v_5489_0;
      if (v_5493_0 == 1) v_5492_0 <= v_5496_0;
      if (v_5500_0 == 1) v_5499_0 <= v_5503_0;
      if (v_5507_0 == 1) v_5506_0 <= v_5510_0;
      if (v_5514_0 == 1) v_5513_0 <= v_5517_0;
      if (v_5521_0 == 1) v_5520_0 <= v_5524_0;
      if (v_5528_0 == 1) v_5527_0 <= v_5531_0;
      if (v_5535_0 == 1) v_5534_0 <= v_5538_0;
      if (v_5542_0 == 1) v_5541_0 <= v_5545_0;
      if (v_5549_0 == 1) v_5548_0 <= v_5552_0;
      if (v_5556_0 == 1) v_5555_0 <= v_5559_0;
      if (v_5563_0 == 1) v_5562_0 <= v_5566_0;
      if (v_5570_0 == 1) v_5569_0 <= v_5573_0;
      if (v_5577_0 == 1) v_5576_0 <= v_5580_0;
      if (v_5584_0 == 1) v_5583_0 <= v_5587_0;
      if (v_5591_0 == 1) v_5590_0 <= v_5594_0;
      if (v_5598_0 == 1) v_5597_0 <= v_5601_0;
      if (v_5605_0 == 1) v_5604_0 <= v_5608_0;
      if (v_5612_0 == 1) v_5611_0 <= v_5615_0;
      if (v_5619_0 == 1) v_5618_0 <= v_5622_0;
      if (v_5626_0 == 1) v_5625_0 <= v_5629_0;
      if (v_5633_0 == 1) v_5632_0 <= v_5636_0;
      if (v_5640_0 == 1) v_5639_0 <= v_5643_0;
      if (v_5647_0 == 1) v_5646_0 <= v_5650_0;
      if (v_5654_0 == 1) v_5653_0 <= v_5657_0;
      if (v_5661_0 == 1) v_5660_0 <= v_5664_0;
      if (v_5668_0 == 1) v_5667_0 <= v_5671_0;
      if (v_5675_0 == 1) v_5674_0 <= v_5678_0;
      if (v_5682_0 == 1) v_5681_0 <= v_5685_0;
      if (v_5689_0 == 1) v_5688_0 <= v_5692_0;
      if (v_5696_0 == 1) v_5695_0 <= v_5699_0;
      if (v_5703_0 == 1) v_5702_0 <= v_5706_0;
      if (v_5710_0 == 1) v_5709_0 <= v_5713_0;
      if (v_5717_0 == 1) v_5716_0 <= v_5720_0;
      if (v_5724_0 == 1) v_5723_0 <= v_5727_0;
      if (v_5731_0 == 1) v_5730_0 <= v_5734_0;
      if (v_5738_0 == 1) v_5737_0 <= v_5741_0;
      if (v_5745_0 == 1) v_5744_0 <= v_5748_0;
      if (v_5752_0 == 1) v_5751_0 <= v_5755_0;
      if (v_5759_0 == 1) v_5758_0 <= v_5762_0;
      if (v_5766_0 == 1) v_5765_0 <= v_5769_0;
      if (v_5773_0 == 1) v_5772_0 <= v_5776_0;
      if (v_5780_0 == 1) v_5779_0 <= v_5783_0;
      if (v_5787_0 == 1) v_5786_0 <= v_5790_0;
      if (v_5794_0 == 1) v_5793_0 <= v_5797_0;
      if (v_5801_0 == 1) v_5800_0 <= v_5804_0;
      if (v_5808_0 == 1) v_5807_0 <= v_5811_0;
      if (v_5815_0 == 1) v_5814_0 <= v_5818_0;
      if (v_5822_0 == 1) v_5821_0 <= v_5825_0;
      if (v_5829_0 == 1) v_5828_0 <= v_5832_0;
      if (v_5836_0 == 1) v_5835_0 <= v_5839_0;
      if (v_5843_0 == 1) v_5842_0 <= v_5846_0;
      if (v_5850_0 == 1) v_5849_0 <= v_5853_0;
      if (v_5857_0 == 1) v_5856_0 <= v_5860_0;
      if (v_5864_0 == 1) v_5863_0 <= v_5867_0;
      if (v_5871_0 == 1) v_5870_0 <= v_5874_0;
      if (v_5878_0 == 1) v_5877_0 <= v_5881_0;
      if (v_5885_0 == 1) v_5884_0 <= v_5888_0;
      if (v_5892_0 == 1) v_5891_0 <= v_5895_0;
      if (v_5899_0 == 1) v_5898_0 <= v_5902_0;
      if (v_5906_0 == 1) v_5905_0 <= v_5909_0;
      if (v_5913_0 == 1) v_5912_0 <= v_5916_0;
      if (v_5920_0 == 1) v_5919_0 <= v_5923_0;
      if (v_5927_0 == 1) v_5926_0 <= v_5930_0;
      if (v_5934_0 == 1) v_5933_0 <= v_5937_0;
      if (v_5941_0 == 1) v_5940_0 <= v_5944_0;
      if (v_5948_0 == 1) v_5947_0 <= v_5951_0;
      if (v_5955_0 == 1) v_5954_0 <= v_5958_0;
      if (v_5962_0 == 1) v_5961_0 <= v_5965_0;
      if (v_5969_0 == 1) v_5968_0 <= v_5972_0;
      if (v_5976_0 == 1) v_5975_0 <= v_5979_0;
      if (v_5983_0 == 1) v_5982_0 <= v_5986_0;
      if (v_5990_0 == 1) v_5989_0 <= v_5993_0;
      if (v_5997_0 == 1) v_5996_0 <= v_6000_0;
      if (v_6004_0 == 1) v_6003_0 <= v_6007_0;
      if (v_6011_0 == 1) v_6010_0 <= v_6014_0;
      if (v_6018_0 == 1) v_6017_0 <= v_6021_0;
      if (v_6025_0 == 1) v_6024_0 <= v_6028_0;
      if (v_6032_0 == 1) v_6031_0 <= v_6035_0;
      if (v_6039_0 == 1) v_6038_0 <= v_6042_0;
      if (v_6046_0 == 1) v_6045_0 <= v_6049_0;
      if (v_6053_0 == 1) v_6052_0 <= v_6056_0;
      if (v_6060_0 == 1) v_6059_0 <= v_6063_0;
      if (v_6067_0 == 1) v_6066_0 <= v_6070_0;
      if (v_6074_0 == 1) v_6073_0 <= v_6077_0;
      if (v_6081_0 == 1) v_6080_0 <= v_6084_0;
      if (v_6088_0 == 1) v_6087_0 <= v_6091_0;
      if (v_6095_0 == 1) v_6094_0 <= v_6098_0;
      if (v_6102_0 == 1) v_6101_0 <= v_6105_0;
      if (v_6109_0 == 1) v_6108_0 <= v_6112_0;
      if (v_6116_0 == 1) v_6115_0 <= v_6119_0;
      if (v_6123_0 == 1) v_6122_0 <= v_6126_0;
      if (v_6130_0 == 1) v_6129_0 <= v_6133_0;
      if (v_6137_0 == 1) v_6136_0 <= v_6140_0;
      if (v_6144_0 == 1) v_6143_0 <= v_6147_0;
      if (v_6151_0 == 1) v_6150_0 <= v_6154_0;
      if (v_6158_0 == 1) v_6157_0 <= v_6161_0;
      if (v_6165_0 == 1) v_6164_0 <= v_6168_0;
      if (v_6172_0 == 1) v_6171_0 <= v_6175_0;
      if (v_6179_0 == 1) v_6178_0 <= v_6182_0;
      if (v_6186_0 == 1) v_6185_0 <= v_6189_0;
      if (v_6193_0 == 1) v_6192_0 <= v_6196_0;
      if (v_6200_0 == 1) v_6199_0 <= v_6203_0;
      if (v_6207_0 == 1) v_6206_0 <= v_6210_0;
      if (v_6214_0 == 1) v_6213_0 <= v_6217_0;
      if (v_6221_0 == 1) v_6220_0 <= v_6224_0;
      if (v_6228_0 == 1) v_6227_0 <= v_6231_0;
      if (v_6235_0 == 1) v_6234_0 <= v_6238_0;
      if (v_6242_0 == 1) v_6241_0 <= v_6245_0;
      if (v_6249_0 == 1) v_6248_0 <= v_6252_0;
      if (v_6256_0 == 1) v_6255_0 <= v_6259_0;
      if (v_6263_0 == 1) v_6262_0 <= v_6266_0;
      if (v_6270_0 == 1) v_6269_0 <= v_6273_0;
      if (v_6277_0 == 1) v_6276_0 <= v_6280_0;
      if (v_6284_0 == 1) v_6283_0 <= v_6287_0;
      if (v_6291_0 == 1) v_6290_0 <= v_6294_0;
      if (v_6298_0 == 1) v_6297_0 <= v_6301_0;
      if (v_6305_0 == 1) v_6304_0 <= v_6308_0;
      if (v_6312_0 == 1) v_6311_0 <= v_6315_0;
      if (v_6319_0 == 1) v_6318_0 <= v_6322_0;
      if (v_6326_0 == 1) v_6325_0 <= v_6329_0;
      if (v_6333_0 == 1) v_6332_0 <= v_6336_0;
      if (v_6340_0 == 1) v_6339_0 <= v_6343_0;
      if (v_6347_0 == 1) v_6346_0 <= v_6350_0;
      if (v_6354_0 == 1) v_6353_0 <= v_6357_0;
      if (v_6361_0 == 1) v_6360_0 <= v_6364_0;
      if (v_6368_0 == 1) v_6367_0 <= v_6371_0;
      if (v_6375_0 == 1) v_6374_0 <= v_6378_0;
      if (v_6382_0 == 1) v_6381_0 <= v_6385_0;
      if (v_6389_0 == 1) v_6388_0 <= v_6392_0;
      if (v_6396_0 == 1) v_6395_0 <= v_6399_0;
      if (v_6403_0 == 1) v_6402_0 <= v_6406_0;
      if (v_6410_0 == 1) v_6409_0 <= v_6413_0;
      if (v_6417_0 == 1) v_6416_0 <= v_6420_0;
      if (v_6424_0 == 1) v_6423_0 <= v_6427_0;
      if (v_6431_0 == 1) v_6430_0 <= v_6434_0;
      if (v_6438_0 == 1) v_6437_0 <= v_6441_0;
      if (v_6445_0 == 1) v_6444_0 <= v_6448_0;
      if (v_6452_0 == 1) v_6451_0 <= v_6455_0;
      if (v_6459_0 == 1) v_6458_0 <= v_6462_0;
      if (v_6466_0 == 1) v_6465_0 <= v_6469_0;
      if (v_6473_0 == 1) v_6472_0 <= v_6476_0;
      if (v_6480_0 == 1) v_6479_0 <= v_6483_0;
      if (v_6487_0 == 1) v_6486_0 <= v_6490_0;
      if (v_6494_0 == 1) v_6493_0 <= v_6497_0;
      if (v_6501_0 == 1) v_6500_0 <= v_6504_0;
      if (v_6508_0 == 1) v_6507_0 <= v_6511_0;
      if (v_6515_0 == 1) v_6514_0 <= v_6518_0;
      if (v_6522_0 == 1) v_6521_0 <= v_6525_0;
      if (v_6529_0 == 1) v_6528_0 <= v_6532_0;
      if (v_6536_0 == 1) v_6535_0 <= v_6539_0;
      if (v_6543_0 == 1) v_6542_0 <= v_6546_0;
      if (v_6550_0 == 1) v_6549_0 <= v_6553_0;
      if (v_6557_0 == 1) v_6556_0 <= v_6560_0;
      if (v_6564_0 == 1) v_6563_0 <= v_6567_0;
      if (v_6571_0 == 1) v_6570_0 <= v_6574_0;
      if (v_6578_0 == 1) v_6577_0 <= v_6581_0;
      if (v_6585_0 == 1) v_6584_0 <= v_6588_0;
      if (v_6592_0 == 1) v_6591_0 <= v_6595_0;
      if (v_6599_0 == 1) v_6598_0 <= v_6602_0;
      if (v_6606_0 == 1) v_6605_0 <= v_6609_0;
      if (v_6613_0 == 1) v_6612_0 <= v_6616_0;
      if (v_6620_0 == 1) v_6619_0 <= v_6623_0;
      if (v_6627_0 == 1) v_6626_0 <= v_6630_0;
      if (v_6634_0 == 1) v_6633_0 <= v_6637_0;
      if (v_6641_0 == 1) v_6640_0 <= v_6644_0;
      if (v_6648_0 == 1) v_6647_0 <= v_6651_0;
      if (v_6655_0 == 1) v_6654_0 <= v_6658_0;
      if (v_6662_0 == 1) v_6661_0 <= v_6665_0;
      if (v_6669_0 == 1) v_6668_0 <= v_6672_0;
      if (v_6676_0 == 1) v_6675_0 <= v_6679_0;
      if (v_6683_0 == 1) v_6682_0 <= v_6686_0;
      if (v_6690_0 == 1) v_6689_0 <= v_6693_0;
      if (v_6697_0 == 1) v_6696_0 <= v_6700_0;
      if (v_6704_0 == 1) v_6703_0 <= v_6707_0;
      if (v_6711_0 == 1) v_6710_0 <= v_6714_0;
      if (v_6718_0 == 1) v_6717_0 <= v_6721_0;
      if (v_6725_0 == 1) v_6724_0 <= v_6728_0;
      if (v_6732_0 == 1) v_6731_0 <= v_6735_0;
      if (v_6739_0 == 1) v_6738_0 <= v_6742_0;
      if (v_6746_0 == 1) v_6745_0 <= v_6749_0;
      if (v_6753_0 == 1) v_6752_0 <= v_6756_0;
      if (v_6760_0 == 1) v_6759_0 <= v_6763_0;
      if (v_6767_0 == 1) v_6766_0 <= v_6770_0;
      if (v_6774_0 == 1) v_6773_0 <= v_6777_0;
      if (v_6781_0 == 1) v_6780_0 <= v_6784_0;
      if (v_6788_0 == 1) v_6787_0 <= v_6791_0;
      if (v_6795_0 == 1) v_6794_0 <= v_6798_0;
      if (v_6802_0 == 1) v_6801_0 <= v_6805_0;
      if (v_6809_0 == 1) v_6808_0 <= v_6812_0;
      if (v_6816_0 == 1) v_6815_0 <= v_6819_0;
      if (v_6823_0 == 1) v_6822_0 <= v_6826_0;
      if (v_6830_0 == 1) v_6829_0 <= v_6833_0;
      if (v_6837_0 == 1) v_6836_0 <= v_6840_0;
      if (v_6844_0 == 1) v_6843_0 <= v_6847_0;
      if (v_6851_0 == 1) v_6850_0 <= v_6854_0;
      if (v_6858_0 == 1) v_6857_0 <= v_6861_0;
      if (v_6865_0 == 1) v_6864_0 <= v_6868_0;
      if (v_6872_0 == 1) v_6871_0 <= v_6875_0;
      if (v_6879_0 == 1) v_6878_0 <= v_6882_0;
      if (v_6886_0 == 1) v_6885_0 <= v_6889_0;
      if (v_6893_0 == 1) v_6892_0 <= v_6896_0;
      if (v_6900_0 == 1) v_6899_0 <= v_6903_0;
      if (v_6907_0 == 1) v_6906_0 <= v_6910_0;
      if (v_6914_0 == 1) v_6913_0 <= v_6917_0;
      if (v_6921_0 == 1) v_6920_0 <= v_6924_0;
      if (v_6928_0 == 1) v_6927_0 <= v_6931_0;
      if (v_6935_0 == 1) v_6934_0 <= v_6938_0;
      if (v_6942_0 == 1) v_6941_0 <= v_6945_0;
      if (v_6949_0 == 1) v_6948_0 <= v_6952_0;
      if (v_6956_0 == 1) v_6955_0 <= v_6959_0;
      if (v_6963_0 == 1) v_6962_0 <= v_6966_0;
      if (v_6970_0 == 1) v_6969_0 <= v_6973_0;
      if (v_6977_0 == 1) v_6976_0 <= v_6980_0;
      if (v_6984_0 == 1) v_6983_0 <= v_6987_0;
      if (v_6991_0 == 1) v_6990_0 <= v_6994_0;
      if (v_6998_0 == 1) v_6997_0 <= v_7001_0;
      if (v_7005_0 == 1) v_7004_0 <= v_7008_0;
      if (v_7012_0 == 1) v_7011_0 <= v_7015_0;
      if (v_7019_0 == 1) v_7018_0 <= v_7022_0;
      if (v_7026_0 == 1) v_7025_0 <= v_7029_0;
      if (v_7033_0 == 1) v_7032_0 <= v_7036_0;
      if (v_7040_0 == 1) v_7039_0 <= v_7043_0;
      if (v_7047_0 == 1) v_7046_0 <= v_7050_0;
      if (v_7054_0 == 1) v_7053_0 <= v_7057_0;
      if (v_7061_0 == 1) v_7060_0 <= v_7064_0;
      if (v_7068_0 == 1) v_7067_0 <= v_7071_0;
      if (v_7075_0 == 1) v_7074_0 <= v_7078_0;
      if (v_7082_0 == 1) v_7081_0 <= v_7085_0;
      if (v_7089_0 == 1) v_7088_0 <= v_7092_0;
      if (v_7096_0 == 1) v_7095_0 <= v_7099_0;
      if (v_7103_0 == 1) v_7102_0 <= v_7106_0;
      if (v_7110_0 == 1) v_7109_0 <= v_7113_0;
      if (v_7117_0 == 1) v_7116_0 <= v_7120_0;
      if (v_7124_0 == 1) v_7123_0 <= v_7127_0;
      if (v_7131_0 == 1) v_7130_0 <= v_7134_0;
      if (v_7138_0 == 1) v_7137_0 <= v_7141_0;
      if (v_7145_0 == 1) v_7144_0 <= v_7148_0;
      if (v_7152_0 == 1) v_7151_0 <= v_7155_0;
      if (v_7159_0 == 1) v_7158_0 <= v_7162_0;
      if (v_7166_0 == 1) v_7165_0 <= v_7169_0;
      if (v_7173_0 == 1) v_7172_0 <= v_7176_0;
      if (v_7180_0 == 1) v_7179_0 <= v_7183_0;
      if (v_7187_0 == 1) v_7186_0 <= v_7190_0;
      if (v_7194_0 == 1) v_7193_0 <= v_7197_0;
      if (v_7201_0 == 1) v_7200_0 <= v_7204_0;
      if (v_7208_0 == 1) v_7207_0 <= v_7211_0;
      if (v_7215_0 == 1) v_7214_0 <= v_7218_0;
      if (v_7222_0 == 1) v_7221_0 <= v_7225_0;
      if (v_7229_0 == 1) v_7228_0 <= v_7232_0;
      if (v_7236_0 == 1) v_7235_0 <= v_7239_0;
      if (v_7243_0 == 1) v_7242_0 <= v_7246_0;
      if (v_7250_0 == 1) v_7249_0 <= v_7253_0;
      if (v_7257_0 == 1) v_7256_0 <= v_7260_0;
      if (v_7264_0 == 1) v_7263_0 <= v_7267_0;
      if (v_7271_0 == 1) v_7270_0 <= v_7274_0;
      if (v_7278_0 == 1) v_7277_0 <= v_7281_0;
      if (v_7285_0 == 1) v_7284_0 <= v_7288_0;
      if (v_7292_0 == 1) v_7291_0 <= v_7295_0;
      if (v_7299_0 == 1) v_7298_0 <= v_7302_0;
      if (v_7306_0 == 1) v_7305_0 <= v_7309_0;
      if (v_7313_0 == 1) v_7312_0 <= v_7316_0;
      if (v_7320_0 == 1) v_7319_0 <= v_7323_0;
      if (v_7327_0 == 1) v_7326_0 <= v_7330_0;
      if (v_7334_0 == 1) v_7333_0 <= v_7337_0;
      if (v_7341_0 == 1) v_7340_0 <= v_7344_0;
      if (v_7348_0 == 1) v_7347_0 <= v_7351_0;
      if (v_7355_0 == 1) v_7354_0 <= v_7358_0;
      if (v_7362_0 == 1) v_7361_0 <= v_7365_0;
      if (v_7369_0 == 1) v_7368_0 <= v_7372_0;
      if (v_7376_0 == 1) v_7375_0 <= v_7379_0;
      if (v_7383_0 == 1) v_7382_0 <= v_7386_0;
      if (v_7390_0 == 1) v_7389_0 <= v_7393_0;
      if (v_7397_0 == 1) v_7396_0 <= v_7400_0;
      if (v_7404_0 == 1) v_7403_0 <= v_7407_0;
      if (v_7411_0 == 1) v_7410_0 <= v_7414_0;
      if (v_7418_0 == 1) v_7417_0 <= v_7421_0;
      if (v_7425_0 == 1) v_7424_0 <= v_7428_0;
      if (v_7432_0 == 1) v_7431_0 <= v_7435_0;
      if (v_7439_0 == 1) v_7438_0 <= v_7442_0;
      if (v_7446_0 == 1) v_7445_0 <= v_7449_0;
      if (v_7453_0 == 1) v_7452_0 <= v_7456_0;
      if (v_7460_0 == 1) v_7459_0 <= v_7463_0;
      if (v_7467_0 == 1) v_7466_0 <= v_7470_0;
      if (v_7474_0 == 1) v_7473_0 <= v_7477_0;
      if (v_7481_0 == 1) v_7480_0 <= v_7484_0;
      if (v_7488_0 == 1) v_7487_0 <= v_7491_0;
      if (v_7495_0 == 1) v_7494_0 <= v_7498_0;
      if (v_7502_0 == 1) v_7501_0 <= v_7505_0;
      if (v_7509_0 == 1) v_7508_0 <= v_7512_0;
      if (v_7516_0 == 1) v_7515_0 <= v_7519_0;
      if (v_7523_0 == 1) v_7522_0 <= v_7526_0;
      if (v_7530_0 == 1) v_7529_0 <= v_7533_0;
      if (v_7537_0 == 1) v_7536_0 <= v_7540_0;
      if (v_7544_0 == 1) v_7543_0 <= v_7547_0;
      if (v_7551_0 == 1) v_7550_0 <= v_7554_0;
      if (v_7558_0 == 1) v_7557_0 <= v_7561_0;
      if (v_7565_0 == 1) v_7564_0 <= v_7568_0;
      if (v_7572_0 == 1) v_7571_0 <= v_7575_0;
      if (v_7579_0 == 1) v_7578_0 <= v_7582_0;
      if (v_7586_0 == 1) v_7585_0 <= v_7589_0;
      if (v_7593_0 == 1) v_7592_0 <= v_7596_0;
      if (v_7600_0 == 1) v_7599_0 <= v_7603_0;
      if (v_7607_0 == 1) v_7606_0 <= v_7610_0;
      if (v_7614_0 == 1) v_7613_0 <= v_7617_0;
      if (v_7621_0 == 1) v_7620_0 <= v_7624_0;
      if (v_7628_0 == 1) v_7627_0 <= v_7631_0;
      if (v_7635_0 == 1) v_7634_0 <= v_7638_0;
      if (v_7642_0 == 1) v_7641_0 <= v_7645_0;
      if (v_7649_0 == 1) v_7648_0 <= v_7652_0;
      if (v_7656_0 == 1) v_7655_0 <= v_7659_0;
      if (v_7663_0 == 1) v_7662_0 <= v_7666_0;
      if (v_7670_0 == 1) v_7669_0 <= v_7673_0;
      if (v_7677_0 == 1) v_7676_0 <= v_7680_0;
      if (v_7684_0 == 1) v_7683_0 <= v_7687_0;
      if (v_7691_0 == 1) v_7690_0 <= v_7694_0;
      if (v_7698_0 == 1) v_7697_0 <= v_7701_0;
      if (v_7705_0 == 1) v_7704_0 <= v_7708_0;
      if (v_7712_0 == 1) v_7711_0 <= v_7715_0;
      if (v_7719_0 == 1) v_7718_0 <= v_7722_0;
      if (v_7726_0 == 1) v_7725_0 <= v_7729_0;
      if (v_7733_0 == 1) v_7732_0 <= v_7736_0;
      if (v_7740_0 == 1) v_7739_0 <= v_7743_0;
      if (v_7747_0 == 1) v_7746_0 <= v_7750_0;
      if (v_7754_0 == 1) v_7753_0 <= v_7757_0;
      if (v_7761_0 == 1) v_7760_0 <= v_7764_0;
      if (v_7768_0 == 1) v_7767_0 <= v_7771_0;
      if (v_7775_0 == 1) v_7774_0 <= v_7778_0;
      if (v_7782_0 == 1) v_7781_0 <= v_7785_0;
      if (v_7789_0 == 1) v_7788_0 <= v_7792_0;
      if (v_7796_0 == 1) v_7795_0 <= v_7799_0;
      if (v_7803_0 == 1) v_7802_0 <= v_7806_0;
      if (v_7810_0 == 1) v_7809_0 <= v_7813_0;
      if (v_7817_0 == 1) v_7816_0 <= v_7820_0;
      if (v_7824_0 == 1) v_7823_0 <= v_7827_0;
      if (v_7831_0 == 1) v_7830_0 <= v_7834_0;
      if (v_7838_0 == 1) v_7837_0 <= v_7841_0;
      if (v_7845_0 == 1) v_7844_0 <= v_7848_0;
      if (v_7852_0 == 1) v_7851_0 <= v_7853_0;
      if (v_11949_0 == 1) v_11948_0 <= v_11954_0;
      v_11960_0 <= 1'h1;
      v_11961_0 <= _act_11962_0;
      v_11965_0 <= v_11966_0;
      if (v_11990_0 == 1) v_11989_0 <= v_11974_0;
      v_11993_0 <= v_11994_0;
      v_12002_0 <= v_12003_0;
      if (v_12066_0 == 1) v_12065_0 <= v_12073_0;
      if (v_12079_0 == 1) v_12078_0 <= v_12080_0;
      if (v_12087_0 == 1) v_12086_0 <= v_12155_0;
      if (v_12087_0 == 1) v_12090_0 <= v_12091_0;
      if (v_12093_0 == 1) v_12092_0 <= v_12143_0;
      if (v_12100_0 == 1) v_12099_0 <= v_12137_0;
      if (1'h1 == 1) v_12109_0 <= v_12103_0;
      if (_act_12111_0 == 1) v_12110_0 <= v_12131_0;
      if (v_12157_0 == 1) v_12156_0 <= v_12165_0;
      v_12170_0 <= 1'h1;
      v_12171_0 <= _act_12111_0;
      v_12173_0 <= v_12174_0;
      v_12178_0 <= v_12179_0;
      v_12183_0 <= v_12184_0;
      if (v_12227_0 == 1) v_12226_0 <= v_12244_0;
      if (v_12268_0 == 1) $write (v_50_0, " ");
      if (v_12270_0 == 1) $write ("    \t[Executed: ", 1'h1, "]", "\n");
      if (v_12272_0 == 1) $write ("Pop", " ");
      if (v_12276_0 == 1) $write
        ("    \t[Executed: ", v_593_0, "]", "\n");
      if (v_12278_0 == 1) $write ("PushPop", " ");
      if (v_12282_0 == 1) $write (v_328_0, " ");
      if (v_12284_0 == 1) $write
        ("    \t[Executed: ", v_628_0, "]", "\n");
      if (v_12286_0 == 1) $write
        ("Impure actions taken (%0d):", v_12289_0, "\n");
      if (v_12286_0 == 1) v_12288_0 <= 1'h1;
      if (v_12292_0 == 1) $finish;
      if (v_14_0 == 1) $write
        ("--All tests passed to depth %0d",
         v_12_0,
         " at time %0d",
         v_12294_0,
         "--",
         "\n");
      if (v_16_0 == 1) v_12294_0 <= v_12295_0;
      if (v_12297_0 == 1) $finish;
      if (v_12299_0 == 1) $write ("Push", " ");
      if (v_12303_0 == 1) $write (v_50_0, " ");
      if (v_12305_0 == 1) $write ("    \t[Executed: ", 1'h1, "]", "\n");
      if (v_12307_0 == 1) $write ("Pop", " ");
      if (v_12311_0 == 1) $write
        ("    \t[Executed: ", v_593_0, "]", "\n");
      if (v_12313_0 == 1) $write ("PushPop", " ");
      if (v_12317_0 == 1) $write (v_328_0, " ");
      if (v_12319_0 == 1) $write
        ("    \t[Executed: ", v_628_0, "]", "\n");
      if (v_19_0 == 1) $write
        ("@ Fail at time %0d", v_12294_0, " @", "\n");
      if (v_12322_0 == 1) $write ("*** ", "StackTopEq", " ");
      if (v_12324_0 == 1) $write ("failed! ***", "\n");
      if (v_12335_0 == 1) v_12334_0 <= v_12344_0;
      if (v_12346_0 == 1) v_12345_0 <= v_12352_0;
      if (v_12335_0 == 1) v_12356_0 <= v_12357_0;
      if (v_12359_0 == 1) v_12358_0 <= v_12367_0;
    end
  end
endmodule