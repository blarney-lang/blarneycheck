// SoC.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module SoC (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         blarneycomponent_0_avalon_master_waitrequest;                // mm_interconnect_0:BlarneyComponent_0_avalon_master_waitrequest -> BlarneyComponent_0:waitrequest
	wire  [31:0] blarneycomponent_0_avalon_master_readdata;                   // mm_interconnect_0:BlarneyComponent_0_avalon_master_readdata -> BlarneyComponent_0:readdata
	wire   [2:0] blarneycomponent_0_avalon_master_address;                    // BlarneyComponent_0:address -> mm_interconnect_0:BlarneyComponent_0_avalon_master_address
	wire         blarneycomponent_0_avalon_master_read;                       // BlarneyComponent_0:read -> mm_interconnect_0:BlarneyComponent_0_avalon_master_read
	wire  [31:0] blarneycomponent_0_avalon_master_writedata;                  // BlarneyComponent_0:writedata -> mm_interconnect_0:BlarneyComponent_0_avalon_master_writedata
	wire         blarneycomponent_0_avalon_master_write;                      // BlarneyComponent_0:write -> mm_interconnect_0:BlarneyComponent_0_avalon_master_write
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [BlarneyComponent_0:reset, jtag_uart_0:rst_n, mm_interconnect_0:BlarneyComponent_0_reset_reset_bridge_in_reset_reset]

	BlarneyComponent blarneycomponent_0 (
		.reset       (rst_controller_reset_out_reset),               //         reset.reset
		.clock       (clk_clk),                                      //         clock.clk
		.address     (blarneycomponent_0_avalon_master_address),     // avalon_master.address
		.writedata   (blarneycomponent_0_avalon_master_writedata),   //              .writedata
		.write       (blarneycomponent_0_avalon_master_write),       //              .write
		.read        (blarneycomponent_0_avalon_master_read),        //              .read
		.waitrequest (blarneycomponent_0_avalon_master_waitrequest), //              .waitrequest
		.readdata    (blarneycomponent_0_avalon_master_readdata)     //              .readdata
	);

	SoC_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         ()                                                             //               irq.irq
	);

	SoC_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                       (clk_clk),                                                     //                                     clk_50_clk.clk
		.BlarneyComponent_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // BlarneyComponent_0_reset_reset_bridge_in_reset.reset
		.BlarneyComponent_0_avalon_master_address             (blarneycomponent_0_avalon_master_address),                    //               BlarneyComponent_0_avalon_master.address
		.BlarneyComponent_0_avalon_master_waitrequest         (blarneycomponent_0_avalon_master_waitrequest),                //                                               .waitrequest
		.BlarneyComponent_0_avalon_master_read                (blarneycomponent_0_avalon_master_read),                       //                                               .read
		.BlarneyComponent_0_avalon_master_readdata            (blarneycomponent_0_avalon_master_readdata),                   //                                               .readdata
		.BlarneyComponent_0_avalon_master_write               (blarneycomponent_0_avalon_master_write),                      //                                               .write
		.BlarneyComponent_0_avalon_master_writedata           (blarneycomponent_0_avalon_master_writedata),                  //                                               .writedata
		.jtag_uart_0_avalon_jtag_slave_address                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                               .write
		.jtag_uart_0_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                               .read
		.jtag_uart_0_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                               .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                               .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                               .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect)   //                                               .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
