module Top
  (input wire clock,
   input wire reset,
   input wire [0:0] in_canPeek,
   input wire [0:0] out_consume_en,
   input wire [7:0] in_peek,
   output wire [0:0] in_consume_en,
   output wire [0:0] out_canPeek,
   output wire [7:0] out_peek);
  // Declarations
  //////////////////////////////////////////////////////////////////////////////
  wire [0:0] v_1_0;
  wire [0:0] v_2_0;
  wire [0:0] v_3_0;
  wire [0:0] v_4_0;
  reg [0:0] v_5_0 = 1'h0;
  wire [0:0] v_6_0;
  wire [0:0] v_7_0;
  wire [0:0] v_8_0;
  wire [0:0] v_9_0;
  wire [0:0] v_10_0;
  wire [0:0] v_11_0;
  reg [0:0] v_12_0 = 1'h0;
  wire [0:0] v_13_0;
  wire [0:0] v_14_0;
  wire [0:0] v_15_0;
  wire [0:0] v_16_0;
  wire [3:0] v_17_0;
  wire [3:0] v_18_0;
  reg [3:0] v_19_0 = 4'h0;
  wire [0:0] v_20_0;
  wire [0:0] v_21_0;
  wire [0:0] v_22_0;
  wire [0:0] v_23_0;
  wire [0:0] v_24_0;
  wire [0:0] v_25_0;
  wire [0:0] v_26_0;
  reg [0:0] v_27_0 = 1'h0;
  wire [0:0] v_28_0;
  wire [0:0] v_29_0;
  wire [0:0] v_30_0;
  wire [0:0] v_31_0;
  wire [0:0] v_32_0;
  wire [0:0] v_33_0;
  wire [0:0] v_34_0;
  wire [0:0] v_35_0;
  wire [0:0] v_36_0;
  wire [0:0] v_37_0;
  reg [3:0] v_38_0 = 4'h0;
  wire [0:0] v_39_0;
  wire [0:0] v_40_0;
  wire [0:0] v_41_0;
  wire [0:0] v_42_0;
  wire [0:0] v_43_0;
  wire [0:0] v_44_0;
  wire [0:0] v_45_0;
  reg [3:0] v_46_0 = 4'h0;
  wire [0:0] v_47_0;
  wire [0:0] v_48_0;
  wire [0:0] v_49_0;
  wire [0:0] v_50_0;
  wire [0:0] v_51_0;
  wire [0:0] v_52_0;
  wire [0:0] v_53_0;
  wire [0:0] v_54_0;
  wire [0:0] v_55_0;
  wire [3:0] v_56_0;
  wire [3:0] v_57_0;
  wire [3:0] v_58_0;
  wire [3:0] v_59_0;
  wire [3:0] v_60_0;
  wire [3:0] v_61_0;
  wire [0:0] v_62_0;
  wire [0:0] v_63_0;
  wire [0:0] v_64_0;
  wire [3:0] v_65_0;
  wire [3:0] v_66_0;
  wire [3:0] v_67_0;
  wire [3:0] v_68_0;
  wire [3:0] v_69_0;
  wire [3:0] v_70_0;
  wire [0:0] v_71_0;
  wire [0:0] v_72_0;
  reg [3:0] v_73_0 = 4'h0;
  wire [0:0] v_74_0;
  wire [0:0] v_75_0;
  wire [0:0] v_76_0;
  wire [0:0] v_77_0;
  wire [0:0] v_78_0;
  wire [0:0] v_79_0;
  wire [0:0] v_80_0;
  reg [3:0] v_81_0 = 4'h0;
  wire [0:0] v_82_0;
  wire [0:0] v_83_0;
  wire [0:0] v_84_0;
  wire [0:0] v_85_0;
  wire [0:0] v_86_0;
  wire [0:0] v_87_0;
  wire [0:0] v_88_0;
  wire [0:0] v_89_0;
  wire [3:0] v_90_0;
  wire [3:0] v_91_0;
  wire [3:0] v_92_0;
  wire [3:0] v_93_0;
  wire [3:0] v_94_0;
  wire [3:0] v_95_0;
  wire [0:0] v_96_0;
  wire [0:0] v_97_0;
  wire [0:0] v_98_0;
  wire [3:0] v_99_0;
  wire [3:0] v_100_0;
  wire [3:0] v_101_0;
  wire [3:0] v_102_0;
  wire [3:0] v_103_0;
  wire [3:0] v_104_0;
  wire [0:0] v_105_0;
  wire [0:0] v_106_0;
  wire [0:0] v_107_0;
  wire [0:0] v_108_0;
  wire [0:0] v_109_0;
  wire [0:0] v_110_0;
  wire [3:0] v_111_0;
  wire [3:0] v_112_0;
  wire [3:0] v_113_0;
  wire [3:0] v_114_0;
  wire [3:0] v_115_0;
  wire [3:0] v_116_0;
  wire [3:0] v_117_0;
  wire [3:0] v_118_0;
  wire [0:0] v_119_0;
  wire [0:0] v_120_0;
  wire [3:0] v_121_0;
  wire [3:0] v_122_0;
  wire [0:0] v_123_0;
  wire [0:0] v_124_0;
  wire [0:0] v_125_0;
  wire [0:0] v_126_0;
  reg [31:0] v_128_0 = 32'h0;
  wire [31:0] v_129_0;
  wire [0:0] v_133_0;
  wire [0:0] v_135_0;
  wire [0:0] v_137_0;
  wire [0:0] v_139_0;
  wire [0:0] v_141_0;
  wire [0:0] v_142_0;
  wire [0:0] v_144_0;
  wire [0:0] v_146_0;
  wire [0:0] v_148_0;
  wire [0:0] v_150_0;
  wire [0:0] v_151_0;
  wire [0:0] v_153_0;
  wire [0:0] v_154_0;
  wire [0:0] v_155_0;
  wire [0:0] v_156_0;
  wire [0:0] v_157_0;
  wire [0:0] v_158_0;
  reg [0:0] v_160_0 = 1'h0;
  wire [0:0] v_161_0;
  wire [0:0] v_162_0;
  wire [0:0] v_163_0;
  wire [0:0] v_164_0;
  wire [0:0] v_165_0;
  wire [0:0] v_166_0;
  wire [0:0] v_167_0;
  wire [0:0] v_168_0;
  wire [0:0] v_169_0;
  wire [0:0] v_170_0;
  reg [0:0] v_171_0 = 1'h0;
  wire [0:0] v_172_0;
  wire [0:0] v_173_0;
  wire [0:0] _act_174_0;
  wire [0:0] v_175_0;
  wire [0:0] v_176_0;
  wire [0:0] v_177_0;
  wire [0:0] v_178_0;
  wire [0:0] v_179_0;
  wire [0:0] v_180_0;
  reg [7:0] v_182_0 = 8'h0;
  wire [7:0] v_183_0;
  reg [7:0] v_184_0 = 8'h0;
  wire [0:0] v_185_0;
  wire [0:0] v_186_0;
  wire [0:0] v_187_0;
  wire [0:0] v_188_0;
  wire [0:0] v_189_0;
  wire [0:0] v_190_0;
  wire [0:0] v_191_0;
  wire [0:0] v_192_0;
  wire [7:0] v_193_0;
  wire [7:0] v_194_0;
  wire [0:0] v_195_0;
  wire [7:0] v_196_0;
  wire [7:0] v_197_0;
  wire [7:0] v_198_0;
  wire [7:0] v_199_0;
  // Instances
  //////////////////////////////////////////////////////////////////////////////
  assign v_1_0 = 1'h1 & v_2_0;
  assign v_2_0 = v_3_0 & v_12_0;
  assign v_3_0 = 1'h1 & v_4_0;
  assign v_4_0 = ~v_5_0;
  assign v_6_0 = v_7_0 | v_1_0;
  assign v_7_0 = v_8_0 & v_123_0;
  assign v_8_0 = v_9_0 & 1'h1;
  assign v_9_0 = v_10_0 & v_25_0;
  assign v_10_0 = v_3_0 & v_11_0;
  assign v_11_0 = ~v_12_0;
  assign v_13_0 = v_14_0 & v_23_0;
  assign v_14_0 = v_15_0 | v_119_0;
  assign v_15_0 = ~v_16_0;
  assign v_16_0 = v_17_0 == v_117_0;
  assign v_17_0 = v_18_0 + v_46_0;
  assign v_18_0 = v_19_0 + v_38_0;
  assign v_20_0 = v_21_0 | v_108_0;
  assign v_21_0 = v_22_0 & v_107_0;
  assign v_22_0 = v_23_0 & v_106_0;
  assign v_23_0 = v_10_0 & v_24_0;
  assign v_24_0 = ~v_25_0;
  assign v_25_0 = v_26_0 | v_27_0;
  assign v_26_0 = ~1'h1;
  assign v_28_0 = v_23_0 | v_29_0;
  assign v_29_0 = v_9_0 & v_30_0;
  assign v_30_0 = ~1'h1;
  assign v_31_0 = v_32_0 | v_105_0;
  assign v_32_0 = v_23_0 ? v_33_0 : 1'h0;
  assign v_33_0 = v_34_0 & v_71_0;
  assign v_34_0 = v_35_0 & v_36_0;
  assign v_35_0 = v_19_0 == 4'hf;
  assign v_36_0 = v_37_0 & v_44_0;
  assign v_37_0 = v_38_0 == 4'hf;
  assign v_39_0 = v_40_0 | v_62_0;
  assign v_40_0 = v_41_0 & v_43_0;
  assign v_41_0 = v_21_0 & v_42_0;
  assign v_42_0 = v_38_0 == 4'hf;
  assign v_43_0 = ~v_44_0;
  assign v_44_0 = v_45_0 & 1'h1;
  assign v_45_0 = v_46_0 == 4'hf;
  assign v_47_0 = v_48_0 | v_52_0;
  assign v_48_0 = v_49_0 & v_51_0;
  assign v_49_0 = v_40_0 & v_50_0;
  assign v_50_0 = v_46_0 == 4'hf;
  assign v_51_0 = ~1'h1;
  assign v_52_0 = v_53_0 | v_54_0;
  assign v_53_0 = v_33_0 & v_23_0;
  assign v_54_0 = v_40_0 & v_55_0;
  assign v_55_0 = ~v_50_0;
  assign v_56_0 = v_57_0 | v_58_0;
  assign v_57_0 = v_48_0 ? 4'h0 : 4'h0;
  assign v_58_0 = v_59_0 | v_60_0;
  assign v_59_0 = v_53_0 ? 4'h0 : 4'h0;
  assign v_60_0 = v_54_0 ? v_61_0 : 4'h0;
  assign v_61_0 = v_46_0 + 4'h1;
  assign v_62_0 = v_53_0 | v_63_0;
  assign v_63_0 = v_21_0 & v_64_0;
  assign v_64_0 = ~v_42_0;
  assign v_65_0 = v_66_0 | v_67_0;
  assign v_66_0 = v_40_0 ? 4'h0 : 4'h0;
  assign v_67_0 = v_68_0 | v_69_0;
  assign v_68_0 = v_53_0 ? 4'h0 : 4'h0;
  assign v_69_0 = v_63_0 ? v_70_0 : 4'h0;
  assign v_70_0 = v_38_0 + 4'h1;
  assign v_71_0 = v_72_0 & v_79_0;
  assign v_72_0 = v_73_0 == 4'hf;
  assign v_74_0 = v_75_0 | v_96_0;
  assign v_75_0 = v_76_0 & v_78_0;
  assign v_76_0 = v_23_0 & v_77_0;
  assign v_77_0 = v_73_0 == 4'hf;
  assign v_78_0 = ~v_79_0;
  assign v_79_0 = v_80_0 & 1'h1;
  assign v_80_0 = v_81_0 == 4'hf;
  assign v_82_0 = v_83_0 | v_87_0;
  assign v_83_0 = v_84_0 & v_86_0;
  assign v_84_0 = v_75_0 & v_85_0;
  assign v_85_0 = v_81_0 == 4'hf;
  assign v_86_0 = ~1'h1;
  assign v_87_0 = v_53_0 | v_88_0;
  assign v_88_0 = v_75_0 & v_89_0;
  assign v_89_0 = ~v_85_0;
  assign v_90_0 = v_91_0 | v_92_0;
  assign v_91_0 = v_83_0 ? 4'h0 : 4'h0;
  assign v_92_0 = v_93_0 | v_94_0;
  assign v_93_0 = v_53_0 ? 4'h0 : 4'h0;
  assign v_94_0 = v_88_0 ? v_95_0 : 4'h0;
  assign v_95_0 = v_81_0 + 4'h1;
  assign v_96_0 = v_53_0 | v_97_0;
  assign v_97_0 = v_23_0 & v_98_0;
  assign v_98_0 = ~v_77_0;
  assign v_99_0 = v_100_0 | v_101_0;
  assign v_100_0 = v_75_0 ? 4'h0 : 4'h0;
  assign v_101_0 = v_102_0 | v_103_0;
  assign v_102_0 = v_53_0 ? 4'h0 : 4'h0;
  assign v_103_0 = v_97_0 ? v_104_0 : 4'h0;
  assign v_104_0 = v_73_0 + 4'h1;
  assign v_105_0 = v_29_0 ? 1'h0 : 1'h0;
  assign v_106_0 = v_19_0 == 4'hf;
  assign v_107_0 = ~v_36_0;
  assign v_108_0 = v_53_0 | v_109_0;
  assign v_109_0 = v_23_0 & v_110_0;
  assign v_110_0 = ~v_106_0;
  assign v_111_0 = v_112_0 | v_113_0;
  assign v_112_0 = v_21_0 ? 4'h0 : 4'h0;
  assign v_113_0 = v_114_0 | v_115_0;
  assign v_114_0 = v_53_0 ? 4'h0 : 4'h0;
  assign v_115_0 = v_109_0 ? v_116_0 : 4'h0;
  assign v_116_0 = v_19_0 + 4'h1;
  assign v_117_0 = v_19_0 + v_118_0;
  assign v_118_0 = v_38_0 + v_46_0;
  assign v_119_0 = ~v_120_0;
  assign v_120_0 = v_121_0 == v_122_0;
  assign v_121_0 = v_73_0 + v_81_0;
  assign v_122_0 = v_81_0 + v_73_0;
  assign v_123_0 = 16'h0 <= 16'h0;
  assign v_124_0 = v_125_0 | v_126_0;
  assign v_125_0 = v_7_0 ? 1'h1 : 1'h0;
  assign v_126_0 = v_1_0 ? 1'h1 : 1'h0;
  assign v_129_0 = v_128_0 + 32'h1;
  assign v_133_0 = v_15_0 & v_13_0;
  assign v_135_0 = v_15_0 & v_13_0;
  assign v_137_0 = v_15_0 & v_13_0;
  assign v_139_0 = v_15_0 & v_13_0;
  assign v_141_0 = v_142_0 & v_13_0;
  assign v_142_0 = ~v_16_0;
  assign v_144_0 = v_119_0 & v_13_0;
  assign v_146_0 = v_119_0 & v_13_0;
  assign v_148_0 = v_119_0 & v_13_0;
  assign v_150_0 = v_151_0 & v_13_0;
  assign v_151_0 = ~v_120_0;
  assign in_consume_en = v_153_0;
  assign v_153_0 = v_154_0 | v_157_0;
  assign v_154_0 = v_155_0 ? 1'h1 : 1'h0;
  assign v_155_0 = v_156_0 & 1'h1;
  assign v_156_0 = in_canPeek;
  assign v_157_0 = v_158_0 ? 1'h0 : 1'h0;
  assign v_158_0 = ~v_155_0;
  assign out_canPeek = v_160_0;
  assign v_161_0 = 1'h1 & v_162_0;
  assign v_162_0 = v_163_0 | v_164_0;
  assign v_163_0 = ~v_160_0;
  assign v_164_0 = v_165_0 | v_168_0;
  assign v_165_0 = v_166_0 ? 1'h1 : 1'h0;
  assign v_166_0 = v_167_0 & 1'h1;
  assign v_167_0 = out_consume_en;
  assign v_168_0 = v_169_0 ? 1'h0 : 1'h0;
  assign v_169_0 = ~v_166_0;
  assign v_170_0 = v_171_0 | _act_174_0;
  assign v_172_0 = v_173_0 | v_177_0;
  assign v_173_0 = _act_174_0 & v_175_0;
  assign _act_174_0 = v_13_0 | v_7_0;
  assign v_175_0 = 1'h1 & v_176_0;
  assign v_176_0 = ~v_162_0;
  assign v_177_0 = v_171_0 & v_161_0;
  assign v_178_0 = v_179_0 | v_180_0;
  assign v_179_0 = v_173_0 ? 1'h1 : 1'h0;
  assign v_180_0 = v_177_0 ? _act_174_0 : 1'h0;
  assign out_peek = v_182_0;
  assign v_183_0 = v_171_0 ? v_184_0 : v_193_0;
  assign v_185_0 = v_186_0 & 1'h1;
  assign v_186_0 = v_187_0 | v_190_0;
  assign v_187_0 = v_188_0 ? 1'h0 : 1'h0;
  assign v_188_0 = ~v_189_0;
  assign v_189_0 = v_173_0 | v_177_0;
  assign v_190_0 = v_191_0 | v_192_0;
  assign v_191_0 = v_173_0 ? 1'h1 : 1'h0;
  assign v_192_0 = v_177_0 ? 1'h1 : 1'h0;
  assign v_193_0 = v_194_0 | v_196_0;
  assign v_194_0 = v_195_0 ? 8'bxxxxxxxx : 8'h0;
  assign v_195_0 = ~_act_174_0;
  assign v_196_0 = v_197_0 | v_198_0;
  assign v_197_0 = v_13_0 ? 8'h46 : 8'h0;
  assign v_198_0 = v_7_0 ? 8'h50 : 8'h0;
  assign v_199_0 = in_peek;
  // Always block
  //////////////////////////////////////////////////////////////////////////////
  always @(posedge clock) begin
    if (reset) begin
      v_5_0 <= 1'h0;
      v_12_0 <= 1'h0;
      v_19_0 <= 4'h0;
      v_27_0 <= 1'h0;
      v_38_0 <= 4'h0;
      v_46_0 <= 4'h0;
      v_73_0 <= 4'h0;
      v_81_0 <= 4'h0;
      v_128_0 <= 32'h0;
      v_160_0 <= 1'h0;
      v_171_0 <= 1'h0;
      v_182_0 <= 8'h0;
      v_184_0 <= 8'h0;
    end else begin
      if (v_1_0 == 1) $finish;
      if (v_6_0 == 1) v_5_0 <= v_124_0;
      if (v_13_0 == 1) v_12_0 <= 1'h1;
      if (v_20_0 == 1) v_19_0 <= v_111_0;
      if (v_28_0 == 1) v_27_0 <= v_31_0;
      if (v_39_0 == 1) v_38_0 <= v_65_0;
      if (v_47_0 == 1) v_46_0 <= v_56_0;
      if (v_74_0 == 1) v_73_0 <= v_99_0;
      if (v_82_0 == 1) v_81_0 <= v_90_0;
      if (v_8_0 == 1) $write
        ("--All tests passed to depth %0d",
         16'h0,
         " at time %0d",
         v_128_0,
         "--",
         "\n");
      if (v_10_0 == 1) v_128_0 <= v_129_0;
      if (v_7_0 == 1) $finish;
      if (v_13_0 == 1) $write
        ("@ Fail at time %0d", v_128_0, " @", "\n");
      if (v_133_0 == 1) $write ("*** ", "Associativity", " ");
      if (v_135_0 == 1) $write (v_19_0, " ");
      if (v_137_0 == 1) $write (v_38_0, " ");
      if (v_139_0 == 1) $write (v_46_0, " ");
      if (v_141_0 == 1) $write ("failed! ***", "\n");
      if (v_144_0 == 1) $write ("*** ", "Commutativity", " ");
      if (v_146_0 == 1) $write (v_73_0, " ");
      if (v_148_0 == 1) $write (v_81_0, " ");
      if (v_150_0 == 1) $write ("failed! ***", "\n");
      if (v_161_0 == 1) v_160_0 <= v_170_0;
      if (v_172_0 == 1) v_171_0 <= v_178_0;
      if (v_161_0 == 1) v_182_0 <= v_183_0;
      if (v_185_0 == 1) v_184_0 <= v_193_0;
    end
  end
endmodule